module main_rt_loopback (
    input  logic        CLOCK_50,
    input  logic [1:0]  KEY,
    input  logic [8:0]  SW,
    input  logic        serial_rx,
    input  logic        dtr_n,
    output logic [6:0]  HEX0,
    output logic [6:0]  HEX1,
    output logic [6:0]  HEX2,
    output logic [6:0]  HEX3,
    output logic [6:0]  HEX4,
    output logic [6:0]  HEX5,
    output logic [7:0]  LED,
    output logic        serial_tx
);

    // === UART RX ===
    logic [7:0] rx_data;
    logic       rx_valid;
    logic [15:0] recv_count;

    uart_rxv2 #(
        .CLK_FREQ(50_000_000),
        .BAUD(115200)
    ) u_rx (
        .clk        (CLOCK_50),
        .rst        (~KEY[0]),
        .serial_rx  (serial_rx),
        .data_out   (rx_data),
        .data_valid (rx_valid),
        .recv_count (recv_count)
    );

    // === UART TX ===
    logic tx_ready;
    logic tx_valid;
    assign tx_valid = rx_valid;   // Direct loopback

    uart_tx #(
        .CLK_FREQ(50_000_000),
        .BAUD(115200)
    ) u_tx (
        .clk        (CLOCK_50),
        .rst        (~KEY[0]),
        .tx_data    (rx_data),
        .tx_valid   (tx_valid),
        .tx_ready   (tx_ready),
        .serial_tx  (serial_tx)
    );

    // === Mode Toggle Logic ===
    logic [2:0] show_mode;
    logic       key1_prev;

    always_ff @(posedge CLOCK_50) begin
        key1_prev <= KEY[1];
        if (~KEY[1] && key1_prev)
            show_mode <= (show_mode == 3) ? 0 : show_mode + 1;
    end

    // === Display Value Selection ===
    logic [23:0] display_val;
    logic [3:0]  mode_val;

    always_comb begin
        case (show_mode)
            3'd0: begin
                display_val = 24'd030314;     // Project ID
                mode_val    = 4'd0;
            end
            3'd1: begin
                display_val = {16'd0, recv_count}; // RX count
                mode_val    = 4'd1;
            end
            3'd2: begin
                display_val = {16'd0, rx_data};    // Latest received
                mode_val    = 4'd2;
            end
            default: begin
                display_val = 24'd999999;
                mode_val    = 4'd0;
            end
        endcase
    end

    // === HEX Display ===
    logic [3:0] digit0, digit1, digit2, digit3, digit4, digit5;

    hex_display u_disp (
        .bin(display_val),
        .digit5(digit5),
        .digit4(digit4),
        .digit3(digit3),
        .digit2(digit2),
        .digit1(digit1),
        .digit0(digit0)
    );

    hex_decoder h0 (.bin(digit0), .seg(HEX0));
    hex_decoder h1 (.bin(digit1), .seg(HEX1));
    hex_decoder h2 (.bin(digit2), .seg(HEX2));
    hex_decoder h3 (.bin(digit3), .seg(HEX3));
    hex_decoder h4 (.bin(digit4), .seg(HEX4));
    hex_decoder h5 (.bin(mode_val), .seg(HEX5));

    // === LED Debugging ===
    assign LED[0] = rx_valid;
    assign LED[1] = tx_valid;
    assign LED[2] = tx_ready;
    assign LED[7:3] = 5'b0;

endmodule
