// fm_wave_gen.sv
module fm_wave_gen1u (
  input  logic        clk,       // your 50 MHz clock
  input  logic        rst,     
  input  logic        in_valid,  // pulse when new rx_data sample is ready
  input  logic [7:0]  in_data,   // filtered sine sample 0–255
  output logic [7:0]  out_data   // FM-modulated sine 0–255
);

  //——— LUT memories —————————————————————————————
  logic [7:0] SINE_LUT [0:1756];
  logic [7:0] STEP_LUT [0:255];

initial begin
    STEP_LUT[0]  = 8'd15;
    STEP_LUT[1]  = 8'd15;
    STEP_LUT[2]  = 8'd15;
    STEP_LUT[3]  = 8'd15;
    STEP_LUT[4]  = 8'd16;
    STEP_LUT[5]  = 8'd16;
    STEP_LUT[6]  = 8'd16;
    STEP_LUT[7]  = 8'd16;
    STEP_LUT[8]  = 8'd16;
    STEP_LUT[9]  = 8'd16;
    STEP_LUT[10]  = 8'd17;
    STEP_LUT[11]  = 8'd17;
    STEP_LUT[12]  = 8'd17;
    STEP_LUT[13]  = 8'd17;
    STEP_LUT[14]  = 8'd17;
    STEP_LUT[15]  = 8'd17;
    STEP_LUT[16]  = 8'd18;
    STEP_LUT[17]  = 8'd18;
    STEP_LUT[18]  = 8'd18;
    STEP_LUT[19]  = 8'd18;
    STEP_LUT[20]  = 8'd18;
    STEP_LUT[21]  = 8'd18;
    STEP_LUT[22]  = 8'd18;
    STEP_LUT[23]  = 8'd19;
    STEP_LUT[24]  = 8'd19;
    STEP_LUT[25]  = 8'd19;
    STEP_LUT[26]  = 8'd19;
    STEP_LUT[27]  = 8'd19;
    STEP_LUT[28]  = 8'd19;
    STEP_LUT[29]  = 8'd20;
    STEP_LUT[30]  = 8'd20;
    STEP_LUT[31]  = 8'd20;
    STEP_LUT[32]  = 8'd20;
    STEP_LUT[33]  = 8'd20;
    STEP_LUT[34]  = 8'd20;
    STEP_LUT[35]  = 8'd20;
    STEP_LUT[36]  = 8'd21;
    STEP_LUT[37]  = 8'd21;
    STEP_LUT[38]  = 8'd21;
    STEP_LUT[39]  = 8'd21;
    STEP_LUT[40]  = 8'd21;
    STEP_LUT[41]  = 8'd21;
    STEP_LUT[42]  = 8'd22;
    STEP_LUT[43]  = 8'd22;
    STEP_LUT[44]  = 8'd22;
    STEP_LUT[45]  = 8'd22;
    STEP_LUT[46]  = 8'd22;
    STEP_LUT[47]  = 8'd22;
    STEP_LUT[48]  = 8'd23;
    STEP_LUT[49]  = 8'd23;
    STEP_LUT[50]  = 8'd23;
    STEP_LUT[51]  = 8'd23;
    STEP_LUT[52]  = 8'd23;
    STEP_LUT[53]  = 8'd23;
    STEP_LUT[54]  = 8'd23;
    STEP_LUT[55]  = 8'd24;
    STEP_LUT[56]  = 8'd24;
    STEP_LUT[57]  = 8'd24;
    STEP_LUT[58]  = 8'd24;
    STEP_LUT[59]  = 8'd24;
    STEP_LUT[60]  = 8'd24;
    STEP_LUT[61]  = 8'd25;
    STEP_LUT[62]  = 8'd25;
    STEP_LUT[63]  = 8'd25;
    STEP_LUT[64]  = 8'd25;
    STEP_LUT[65]  = 8'd25;
    STEP_LUT[66]  = 8'd25;
    STEP_LUT[67]  = 8'd26;
    STEP_LUT[68]  = 8'd26;
    STEP_LUT[69]  = 8'd26;
    STEP_LUT[70]  = 8'd26;
    STEP_LUT[71]  = 8'd26;
    STEP_LUT[72]  = 8'd26;
    STEP_LUT[73]  = 8'd26;
    STEP_LUT[74]  = 8'd27;
    STEP_LUT[75]  = 8'd27;
    STEP_LUT[76]  = 8'd27;
    STEP_LUT[77]  = 8'd27;
    STEP_LUT[78]  = 8'd27;
    STEP_LUT[79]  = 8'd27;
    STEP_LUT[80]  = 8'd28;
    STEP_LUT[81]  = 8'd28;
    STEP_LUT[82]  = 8'd28;
    STEP_LUT[83]  = 8'd28;
    STEP_LUT[84]  = 8'd28;
    STEP_LUT[85]  = 8'd28;
    STEP_LUT[86]  = 8'd28;
    STEP_LUT[87]  = 8'd29;
    STEP_LUT[88]  = 8'd29;
    STEP_LUT[89]  = 8'd29;
    STEP_LUT[90]  = 8'd29;
    STEP_LUT[91]  = 8'd29;
    STEP_LUT[92]  = 8'd29;
    STEP_LUT[93]  = 8'd30;
    STEP_LUT[94]  = 8'd30;
    STEP_LUT[95]  = 8'd30;
    STEP_LUT[96]  = 8'd30;
    STEP_LUT[97]  = 8'd30;
    STEP_LUT[98]  = 8'd30;
    STEP_LUT[99]  = 8'd31;
    STEP_LUT[100]  = 8'd31;
    STEP_LUT[101]  = 8'd31;
    STEP_LUT[102]  = 8'd31;
    STEP_LUT[103]  = 8'd31;
    STEP_LUT[104]  = 8'd31;
    STEP_LUT[105]  = 8'd31;
    STEP_LUT[106]  = 8'd32;
    STEP_LUT[107]  = 8'd32;
    STEP_LUT[108]  = 8'd32;
    STEP_LUT[109]  = 8'd32;
    STEP_LUT[110]  = 8'd32;
    STEP_LUT[111]  = 8'd32;
    STEP_LUT[112]  = 8'd33;
    STEP_LUT[113]  = 8'd33;
    STEP_LUT[114]  = 8'd33;
    STEP_LUT[115]  = 8'd33;
    STEP_LUT[116]  = 8'd33;
    STEP_LUT[117]  = 8'd33;
    STEP_LUT[118]  = 8'd34;
    STEP_LUT[119]  = 8'd34;
    STEP_LUT[120]  = 8'd34;
    STEP_LUT[121]  = 8'd34;
    STEP_LUT[122]  = 8'd34;
    STEP_LUT[123]  = 8'd34;
    STEP_LUT[124]  = 8'd34;
    STEP_LUT[125]  = 8'd35;
    STEP_LUT[126]  = 8'd35;
    STEP_LUT[127]  = 8'd35;
    STEP_LUT[128]  = 8'd35;
    STEP_LUT[129]  = 8'd35;
    STEP_LUT[130]  = 8'd35;
    STEP_LUT[131]  = 8'd36;
    STEP_LUT[132]  = 8'd36;
    STEP_LUT[133]  = 8'd36;
    STEP_LUT[134]  = 8'd36;
    STEP_LUT[135]  = 8'd36;
    STEP_LUT[136]  = 8'd36;
    STEP_LUT[137]  = 8'd36;
    STEP_LUT[138]  = 8'd37;
    STEP_LUT[139]  = 8'd37;
    STEP_LUT[140]  = 8'd37;
    STEP_LUT[141]  = 8'd37;
    STEP_LUT[142]  = 8'd37;
    STEP_LUT[143]  = 8'd37;
    STEP_LUT[144]  = 8'd38;
    STEP_LUT[145]  = 8'd38;
    STEP_LUT[146]  = 8'd38;
    STEP_LUT[147]  = 8'd38;
    STEP_LUT[148]  = 8'd38;
    STEP_LUT[149]  = 8'd38;
    STEP_LUT[150]  = 8'd39;
    STEP_LUT[151]  = 8'd39;
    STEP_LUT[152]  = 8'd39;
    STEP_LUT[153]  = 8'd39;
    STEP_LUT[154]  = 8'd39;
    STEP_LUT[155]  = 8'd39;
    STEP_LUT[156]  = 8'd39;
    STEP_LUT[157]  = 8'd40;
    STEP_LUT[158]  = 8'd40;
    STEP_LUT[159]  = 8'd40;
    STEP_LUT[160]  = 8'd40;
    STEP_LUT[161]  = 8'd40;
    STEP_LUT[162]  = 8'd40;
    STEP_LUT[163]  = 8'd41;
    STEP_LUT[164]  = 8'd41;
    STEP_LUT[165]  = 8'd41;
    STEP_LUT[166]  = 8'd41;
    STEP_LUT[167]  = 8'd41;
    STEP_LUT[168]  = 8'd41;
    STEP_LUT[169]  = 8'd42;
    STEP_LUT[170]  = 8'd42;
    STEP_LUT[171]  = 8'd42;
    STEP_LUT[172]  = 8'd42;
    STEP_LUT[173]  = 8'd42;
    STEP_LUT[174]  = 8'd42;
    STEP_LUT[175]  = 8'd42;
    STEP_LUT[176]  = 8'd43;
    STEP_LUT[177]  = 8'd43;
    STEP_LUT[178]  = 8'd43;
    STEP_LUT[179]  = 8'd43;
    STEP_LUT[180]  = 8'd43;
    STEP_LUT[181]  = 8'd43;
    STEP_LUT[182]  = 8'd44;
    STEP_LUT[183]  = 8'd44;
    STEP_LUT[184]  = 8'd44;
    STEP_LUT[185]  = 8'd44;
    STEP_LUT[186]  = 8'd44;
    STEP_LUT[187]  = 8'd44;
    STEP_LUT[188]  = 8'd44;
    STEP_LUT[189]  = 8'd45;
    STEP_LUT[190]  = 8'd45;
    STEP_LUT[191]  = 8'd45;
    STEP_LUT[192]  = 8'd45;
    STEP_LUT[193]  = 8'd45;
    STEP_LUT[194]  = 8'd45;
    STEP_LUT[195]  = 8'd46;
    STEP_LUT[196]  = 8'd46;
    STEP_LUT[197]  = 8'd46;
    STEP_LUT[198]  = 8'd46;
    STEP_LUT[199]  = 8'd46;
    STEP_LUT[200]  = 8'd46;
    STEP_LUT[201]  = 8'd47;
    STEP_LUT[202]  = 8'd47;
    STEP_LUT[203]  = 8'd47;
    STEP_LUT[204]  = 8'd47;
    STEP_LUT[205]  = 8'd47;
    STEP_LUT[206]  = 8'd47;
    STEP_LUT[207]  = 8'd47;
    STEP_LUT[208]  = 8'd48;
    STEP_LUT[209]  = 8'd48;
    STEP_LUT[210]  = 8'd48;
    STEP_LUT[211]  = 8'd48;
    STEP_LUT[212]  = 8'd48;
    STEP_LUT[213]  = 8'd48;
    STEP_LUT[214]  = 8'd49;
    STEP_LUT[215]  = 8'd49;
    STEP_LUT[216]  = 8'd49;
    STEP_LUT[217]  = 8'd49;
    STEP_LUT[218]  = 8'd49;
    STEP_LUT[219]  = 8'd49;
    STEP_LUT[220]  = 8'd50;
    STEP_LUT[221]  = 8'd50;
    STEP_LUT[222]  = 8'd50;
    STEP_LUT[223]  = 8'd50;
    STEP_LUT[224]  = 8'd50;
    STEP_LUT[225]  = 8'd50;
    STEP_LUT[226]  = 8'd50;
    STEP_LUT[227]  = 8'd51;
    STEP_LUT[228]  = 8'd51;
    STEP_LUT[229]  = 8'd51;
    STEP_LUT[230]  = 8'd51;
    STEP_LUT[231]  = 8'd51;
    STEP_LUT[232]  = 8'd51;
    STEP_LUT[233]  = 8'd52;
    STEP_LUT[234]  = 8'd52;
    STEP_LUT[235]  = 8'd52;
    STEP_LUT[236]  = 8'd52;
    STEP_LUT[237]  = 8'd52;
    STEP_LUT[238]  = 8'd52;
    STEP_LUT[239]  = 8'd52;
    STEP_LUT[240]  = 8'd53;
    STEP_LUT[241]  = 8'd53;
    STEP_LUT[242]  = 8'd53;
    STEP_LUT[243]  = 8'd53;
    STEP_LUT[244]  = 8'd53;
    STEP_LUT[245]  = 8'd53;
    STEP_LUT[246]  = 8'd54;
    STEP_LUT[247]  = 8'd54;
    STEP_LUT[248]  = 8'd54;
    STEP_LUT[249]  = 8'd54;
    STEP_LUT[250]  = 8'd54;
    STEP_LUT[251]  = 8'd54;
    STEP_LUT[252]  = 8'd55;
    STEP_LUT[253]  = 8'd55;
    STEP_LUT[254]  = 8'd55;
    STEP_LUT[255]  = 8'd55;
end


initial begin
    SINE_LUT[0]  = 8'd128;
    SINE_LUT[1]  = 8'd128;
    SINE_LUT[2]  = 8'd129;
    SINE_LUT[3]  = 8'd129;
    SINE_LUT[4]  = 8'd130;
    SINE_LUT[5]  = 8'd130;
    SINE_LUT[6]  = 8'd131;
    SINE_LUT[7]  = 8'd131;
    SINE_LUT[8]  = 8'd132;
    SINE_LUT[9]  = 8'd132;
    SINE_LUT[10]  = 8'd133;
    SINE_LUT[11]  = 8'd133;
    SINE_LUT[12]  = 8'd133;
    SINE_LUT[13]  = 8'd134;
    SINE_LUT[14]  = 8'd134;
    SINE_LUT[15]  = 8'd135;
    SINE_LUT[16]  = 8'd135;
    SINE_LUT[17]  = 8'd136;
    SINE_LUT[18]  = 8'd136;
    SINE_LUT[19]  = 8'd137;
    SINE_LUT[20]  = 8'd137;
    SINE_LUT[21]  = 8'd138;
    SINE_LUT[22]  = 8'd138;
    SINE_LUT[23]  = 8'd138;
    SINE_LUT[24]  = 8'd139;
    SINE_LUT[25]  = 8'd139;
    SINE_LUT[26]  = 8'd140;
    SINE_LUT[27]  = 8'd140;
    SINE_LUT[28]  = 8'd141;
    SINE_LUT[29]  = 8'd141;
    SINE_LUT[30]  = 8'd142;
    SINE_LUT[31]  = 8'd142;
    SINE_LUT[32]  = 8'd143;
    SINE_LUT[33]  = 8'd143;
    SINE_LUT[34]  = 8'd143;
    SINE_LUT[35]  = 8'd144;
    SINE_LUT[36]  = 8'd144;
    SINE_LUT[37]  = 8'd145;
    SINE_LUT[38]  = 8'd145;
    SINE_LUT[39]  = 8'd146;
    SINE_LUT[40]  = 8'd146;
    SINE_LUT[41]  = 8'd147;
    SINE_LUT[42]  = 8'd147;
    SINE_LUT[43]  = 8'd147;
    SINE_LUT[44]  = 8'd148;
    SINE_LUT[45]  = 8'd148;
    SINE_LUT[46]  = 8'd149;
    SINE_LUT[47]  = 8'd149;
    SINE_LUT[48]  = 8'd150;
    SINE_LUT[49]  = 8'd150;
    SINE_LUT[50]  = 8'd151;
    SINE_LUT[51]  = 8'd151;
    SINE_LUT[52]  = 8'd151;
    SINE_LUT[53]  = 8'd152;
    SINE_LUT[54]  = 8'd152;
    SINE_LUT[55]  = 8'd153;
    SINE_LUT[56]  = 8'd153;
    SINE_LUT[57]  = 8'd154;
    SINE_LUT[58]  = 8'd154;
    SINE_LUT[59]  = 8'd155;
    SINE_LUT[60]  = 8'd155;
    SINE_LUT[61]  = 8'd155;
    SINE_LUT[62]  = 8'd156;
    SINE_LUT[63]  = 8'd156;
    SINE_LUT[64]  = 8'd157;
    SINE_LUT[65]  = 8'd157;
    SINE_LUT[66]  = 8'd158;
    SINE_LUT[67]  = 8'd158;
    SINE_LUT[68]  = 8'd159;
    SINE_LUT[69]  = 8'd159;
    SINE_LUT[70]  = 8'd159;
    SINE_LUT[71]  = 8'd160;
    SINE_LUT[72]  = 8'd160;
    SINE_LUT[73]  = 8'd161;
    SINE_LUT[74]  = 8'd161;
    SINE_LUT[75]  = 8'd162;
    SINE_LUT[76]  = 8'd162;
    SINE_LUT[77]  = 8'd163;
    SINE_LUT[78]  = 8'd163;
    SINE_LUT[79]  = 8'd163;
    SINE_LUT[80]  = 8'd164;
    SINE_LUT[81]  = 8'd164;
    SINE_LUT[82]  = 8'd165;
    SINE_LUT[83]  = 8'd165;
    SINE_LUT[84]  = 8'd166;
    SINE_LUT[85]  = 8'd166;
    SINE_LUT[86]  = 8'd166;
    SINE_LUT[87]  = 8'd167;
    SINE_LUT[88]  = 8'd167;
    SINE_LUT[89]  = 8'd168;
    SINE_LUT[90]  = 8'd168;
    SINE_LUT[91]  = 8'd169;
    SINE_LUT[92]  = 8'd169;
    SINE_LUT[93]  = 8'd169;
    SINE_LUT[94]  = 8'd170;
    SINE_LUT[95]  = 8'd170;
    SINE_LUT[96]  = 8'd171;
    SINE_LUT[97]  = 8'd171;
    SINE_LUT[98]  = 8'd172;
    SINE_LUT[99]  = 8'd172;
    SINE_LUT[100]  = 8'd172;
    SINE_LUT[101]  = 8'd173;
    SINE_LUT[102]  = 8'd173;
    SINE_LUT[103]  = 8'd174;
    SINE_LUT[104]  = 8'd174;
    SINE_LUT[105]  = 8'd175;
    SINE_LUT[106]  = 8'd175;
    SINE_LUT[107]  = 8'd175;
    SINE_LUT[108]  = 8'd176;
    SINE_LUT[109]  = 8'd176;
    SINE_LUT[110]  = 8'd177;
    SINE_LUT[111]  = 8'd177;
    SINE_LUT[112]  = 8'd178;
    SINE_LUT[113]  = 8'd178;
    SINE_LUT[114]  = 8'd178;
    SINE_LUT[115]  = 8'd179;
    SINE_LUT[116]  = 8'd179;
    SINE_LUT[117]  = 8'd180;
    SINE_LUT[118]  = 8'd180;
    SINE_LUT[119]  = 8'd180;
    SINE_LUT[120]  = 8'd181;
    SINE_LUT[121]  = 8'd181;
    SINE_LUT[122]  = 8'd182;
    SINE_LUT[123]  = 8'd182;
    SINE_LUT[124]  = 8'd182;
    SINE_LUT[125]  = 8'd183;
    SINE_LUT[126]  = 8'd183;
    SINE_LUT[127]  = 8'd184;
    SINE_LUT[128]  = 8'd184;
    SINE_LUT[129]  = 8'd185;
    SINE_LUT[130]  = 8'd185;
    SINE_LUT[131]  = 8'd185;
    SINE_LUT[132]  = 8'd186;
    SINE_LUT[133]  = 8'd186;
    SINE_LUT[134]  = 8'd187;
    SINE_LUT[135]  = 8'd187;
    SINE_LUT[136]  = 8'd187;
    SINE_LUT[137]  = 8'd188;
    SINE_LUT[138]  = 8'd188;
    SINE_LUT[139]  = 8'd189;
    SINE_LUT[140]  = 8'd189;
    SINE_LUT[141]  = 8'd189;
    SINE_LUT[142]  = 8'd190;
    SINE_LUT[143]  = 8'd190;
    SINE_LUT[144]  = 8'd191;
    SINE_LUT[145]  = 8'd191;
    SINE_LUT[146]  = 8'd191;
    SINE_LUT[147]  = 8'd192;
    SINE_LUT[148]  = 8'd192;
    SINE_LUT[149]  = 8'd193;
    SINE_LUT[150]  = 8'd193;
    SINE_LUT[151]  = 8'd193;
    SINE_LUT[152]  = 8'd194;
    SINE_LUT[153]  = 8'd194;
    SINE_LUT[154]  = 8'd194;
    SINE_LUT[155]  = 8'd195;
    SINE_LUT[156]  = 8'd195;
    SINE_LUT[157]  = 8'd196;
    SINE_LUT[158]  = 8'd196;
    SINE_LUT[159]  = 8'd196;
    SINE_LUT[160]  = 8'd197;
    SINE_LUT[161]  = 8'd197;
    SINE_LUT[162]  = 8'd198;
    SINE_LUT[163]  = 8'd198;
    SINE_LUT[164]  = 8'd198;
    SINE_LUT[165]  = 8'd199;
    SINE_LUT[166]  = 8'd199;
    SINE_LUT[167]  = 8'd199;
    SINE_LUT[168]  = 8'd200;
    SINE_LUT[169]  = 8'd200;
    SINE_LUT[170]  = 8'd201;
    SINE_LUT[171]  = 8'd201;
    SINE_LUT[172]  = 8'd201;
    SINE_LUT[173]  = 8'd202;
    SINE_LUT[174]  = 8'd202;
    SINE_LUT[175]  = 8'd202;
    SINE_LUT[176]  = 8'd203;
    SINE_LUT[177]  = 8'd203;
    SINE_LUT[178]  = 8'd203;
    SINE_LUT[179]  = 8'd204;
    SINE_LUT[180]  = 8'd204;
    SINE_LUT[181]  = 8'd205;
    SINE_LUT[182]  = 8'd205;
    SINE_LUT[183]  = 8'd205;
    SINE_LUT[184]  = 8'd206;
    SINE_LUT[185]  = 8'd206;
    SINE_LUT[186]  = 8'd206;
    SINE_LUT[187]  = 8'd207;
    SINE_LUT[188]  = 8'd207;
    SINE_LUT[189]  = 8'd207;
    SINE_LUT[190]  = 8'd208;
    SINE_LUT[191]  = 8'd208;
    SINE_LUT[192]  = 8'd209;
    SINE_LUT[193]  = 8'd209;
    SINE_LUT[194]  = 8'd209;
    SINE_LUT[195]  = 8'd210;
    SINE_LUT[196]  = 8'd210;
    SINE_LUT[197]  = 8'd210;
    SINE_LUT[198]  = 8'd211;
    SINE_LUT[199]  = 8'd211;
    SINE_LUT[200]  = 8'd211;
    SINE_LUT[201]  = 8'd212;
    SINE_LUT[202]  = 8'd212;
    SINE_LUT[203]  = 8'd212;
    SINE_LUT[204]  = 8'd213;
    SINE_LUT[205]  = 8'd213;
    SINE_LUT[206]  = 8'd213;
    SINE_LUT[207]  = 8'd214;
    SINE_LUT[208]  = 8'd214;
    SINE_LUT[209]  = 8'd214;
    SINE_LUT[210]  = 8'd215;
    SINE_LUT[211]  = 8'd215;
    SINE_LUT[212]  = 8'd215;
    SINE_LUT[213]  = 8'd216;
    SINE_LUT[214]  = 8'd216;
    SINE_LUT[215]  = 8'd216;
    SINE_LUT[216]  = 8'd217;
    SINE_LUT[217]  = 8'd217;
    SINE_LUT[218]  = 8'd217;
    SINE_LUT[219]  = 8'd218;
    SINE_LUT[220]  = 8'd218;
    SINE_LUT[221]  = 8'd218;
    SINE_LUT[222]  = 8'd219;
    SINE_LUT[223]  = 8'd219;
    SINE_LUT[224]  = 8'd219;
    SINE_LUT[225]  = 8'd220;
    SINE_LUT[226]  = 8'd220;
    SINE_LUT[227]  = 8'd220;
    SINE_LUT[228]  = 8'd220;
    SINE_LUT[229]  = 8'd221;
    SINE_LUT[230]  = 8'd221;
    SINE_LUT[231]  = 8'd221;
    SINE_LUT[232]  = 8'd222;
    SINE_LUT[233]  = 8'd222;
    SINE_LUT[234]  = 8'd222;
    SINE_LUT[235]  = 8'd223;
    SINE_LUT[236]  = 8'd223;
    SINE_LUT[237]  = 8'd223;
    SINE_LUT[238]  = 8'd224;
    SINE_LUT[239]  = 8'd224;
    SINE_LUT[240]  = 8'd224;
    SINE_LUT[241]  = 8'd224;
    SINE_LUT[242]  = 8'd225;
    SINE_LUT[243]  = 8'd225;
    SINE_LUT[244]  = 8'd225;
    SINE_LUT[245]  = 8'd226;
    SINE_LUT[246]  = 8'd226;
    SINE_LUT[247]  = 8'd226;
    SINE_LUT[248]  = 8'd226;
    SINE_LUT[249]  = 8'd227;
    SINE_LUT[250]  = 8'd227;
    SINE_LUT[251]  = 8'd227;
    SINE_LUT[252]  = 8'd228;
    SINE_LUT[253]  = 8'd228;
    SINE_LUT[254]  = 8'd228;
    SINE_LUT[255]  = 8'd228;
    SINE_LUT[256]  = 8'd229;
    SINE_LUT[257]  = 8'd229;
    SINE_LUT[258]  = 8'd229;
    SINE_LUT[259]  = 8'd230;
    SINE_LUT[260]  = 8'd230;
    SINE_LUT[261]  = 8'd230;
    SINE_LUT[262]  = 8'd230;
    SINE_LUT[263]  = 8'd231;
    SINE_LUT[264]  = 8'd231;
    SINE_LUT[265]  = 8'd231;
    SINE_LUT[266]  = 8'd231;
    SINE_LUT[267]  = 8'd232;
    SINE_LUT[268]  = 8'd232;
    SINE_LUT[269]  = 8'd232;
    SINE_LUT[270]  = 8'd232;
    SINE_LUT[271]  = 8'd233;
    SINE_LUT[272]  = 8'd233;
    SINE_LUT[273]  = 8'd233;
    SINE_LUT[274]  = 8'd233;
    SINE_LUT[275]  = 8'd234;
    SINE_LUT[276]  = 8'd234;
    SINE_LUT[277]  = 8'd234;
    SINE_LUT[278]  = 8'd234;
    SINE_LUT[279]  = 8'd235;
    SINE_LUT[280]  = 8'd235;
    SINE_LUT[281]  = 8'd235;
    SINE_LUT[282]  = 8'd235;
    SINE_LUT[283]  = 8'd236;
    SINE_LUT[284]  = 8'd236;
    SINE_LUT[285]  = 8'd236;
    SINE_LUT[286]  = 8'd236;
    SINE_LUT[287]  = 8'd237;
    SINE_LUT[288]  = 8'd237;
    SINE_LUT[289]  = 8'd237;
    SINE_LUT[290]  = 8'd237;
    SINE_LUT[291]  = 8'd238;
    SINE_LUT[292]  = 8'd238;
    SINE_LUT[293]  = 8'd238;
    SINE_LUT[294]  = 8'd238;
    SINE_LUT[295]  = 8'd238;
    SINE_LUT[296]  = 8'd239;
    SINE_LUT[297]  = 8'd239;
    SINE_LUT[298]  = 8'd239;
    SINE_LUT[299]  = 8'd239;
    SINE_LUT[300]  = 8'd240;
    SINE_LUT[301]  = 8'd240;
    SINE_LUT[302]  = 8'd240;
    SINE_LUT[303]  = 8'd240;
    SINE_LUT[304]  = 8'd240;
    SINE_LUT[305]  = 8'd241;
    SINE_LUT[306]  = 8'd241;
    SINE_LUT[307]  = 8'd241;
    SINE_LUT[308]  = 8'd241;
    SINE_LUT[309]  = 8'd241;
    SINE_LUT[310]  = 8'd242;
    SINE_LUT[311]  = 8'd242;
    SINE_LUT[312]  = 8'd242;
    SINE_LUT[313]  = 8'd242;
    SINE_LUT[314]  = 8'd242;
    SINE_LUT[315]  = 8'd243;
    SINE_LUT[316]  = 8'd243;
    SINE_LUT[317]  = 8'd243;
    SINE_LUT[318]  = 8'd243;
    SINE_LUT[319]  = 8'd243;
    SINE_LUT[320]  = 8'd244;
    SINE_LUT[321]  = 8'd244;
    SINE_LUT[322]  = 8'd244;
    SINE_LUT[323]  = 8'd244;
    SINE_LUT[324]  = 8'd244;
    SINE_LUT[325]  = 8'd245;
    SINE_LUT[326]  = 8'd245;
    SINE_LUT[327]  = 8'd245;
    SINE_LUT[328]  = 8'd245;
    SINE_LUT[329]  = 8'd245;
    SINE_LUT[330]  = 8'd245;
    SINE_LUT[331]  = 8'd246;
    SINE_LUT[332]  = 8'd246;
    SINE_LUT[333]  = 8'd246;
    SINE_LUT[334]  = 8'd246;
    SINE_LUT[335]  = 8'd246;
    SINE_LUT[336]  = 8'd246;
    SINE_LUT[337]  = 8'd247;
    SINE_LUT[338]  = 8'd247;
    SINE_LUT[339]  = 8'd247;
    SINE_LUT[340]  = 8'd247;
    SINE_LUT[341]  = 8'd247;
    SINE_LUT[342]  = 8'd247;
    SINE_LUT[343]  = 8'd248;
    SINE_LUT[344]  = 8'd248;
    SINE_LUT[345]  = 8'd248;
    SINE_LUT[346]  = 8'd248;
    SINE_LUT[347]  = 8'd248;
    SINE_LUT[348]  = 8'd248;
    SINE_LUT[349]  = 8'd248;
    SINE_LUT[350]  = 8'd249;
    SINE_LUT[351]  = 8'd249;
    SINE_LUT[352]  = 8'd249;
    SINE_LUT[353]  = 8'd249;
    SINE_LUT[354]  = 8'd249;
    SINE_LUT[355]  = 8'd249;
    SINE_LUT[356]  = 8'd249;
    SINE_LUT[357]  = 8'd250;
    SINE_LUT[358]  = 8'd250;
    SINE_LUT[359]  = 8'd250;
    SINE_LUT[360]  = 8'd250;
    SINE_LUT[361]  = 8'd250;
    SINE_LUT[362]  = 8'd250;
    SINE_LUT[363]  = 8'd250;
    SINE_LUT[364]  = 8'd250;
    SINE_LUT[365]  = 8'd251;
    SINE_LUT[366]  = 8'd251;
    SINE_LUT[367]  = 8'd251;
    SINE_LUT[368]  = 8'd251;
    SINE_LUT[369]  = 8'd251;
    SINE_LUT[370]  = 8'd251;
    SINE_LUT[371]  = 8'd251;
    SINE_LUT[372]  = 8'd251;
    SINE_LUT[373]  = 8'd251;
    SINE_LUT[374]  = 8'd252;
    SINE_LUT[375]  = 8'd252;
    SINE_LUT[376]  = 8'd252;
    SINE_LUT[377]  = 8'd252;
    SINE_LUT[378]  = 8'd252;
    SINE_LUT[379]  = 8'd252;
    SINE_LUT[380]  = 8'd252;
    SINE_LUT[381]  = 8'd252;
    SINE_LUT[382]  = 8'd252;
    SINE_LUT[383]  = 8'd252;
    SINE_LUT[384]  = 8'd253;
    SINE_LUT[385]  = 8'd253;
    SINE_LUT[386]  = 8'd253;
    SINE_LUT[387]  = 8'd253;
    SINE_LUT[388]  = 8'd253;
    SINE_LUT[389]  = 8'd253;
    SINE_LUT[390]  = 8'd253;
    SINE_LUT[391]  = 8'd253;
    SINE_LUT[392]  = 8'd253;
    SINE_LUT[393]  = 8'd253;
    SINE_LUT[394]  = 8'd253;
    SINE_LUT[395]  = 8'd253;
    SINE_LUT[396]  = 8'd253;
    SINE_LUT[397]  = 8'd254;
    SINE_LUT[398]  = 8'd254;
    SINE_LUT[399]  = 8'd254;
    SINE_LUT[400]  = 8'd254;
    SINE_LUT[401]  = 8'd254;
    SINE_LUT[402]  = 8'd254;
    SINE_LUT[403]  = 8'd254;
    SINE_LUT[404]  = 8'd254;
    SINE_LUT[405]  = 8'd254;
    SINE_LUT[406]  = 8'd254;
    SINE_LUT[407]  = 8'd254;
    SINE_LUT[408]  = 8'd254;
    SINE_LUT[409]  = 8'd254;
    SINE_LUT[410]  = 8'd254;
    SINE_LUT[411]  = 8'd254;
    SINE_LUT[412]  = 8'd254;
    SINE_LUT[413]  = 8'd254;
    SINE_LUT[414]  = 8'd254;
    SINE_LUT[415]  = 8'd255;
    SINE_LUT[416]  = 8'd255;
    SINE_LUT[417]  = 8'd255;
    SINE_LUT[418]  = 8'd255;
    SINE_LUT[419]  = 8'd255;
    SINE_LUT[420]  = 8'd255;
    SINE_LUT[421]  = 8'd255;
    SINE_LUT[422]  = 8'd255;
    SINE_LUT[423]  = 8'd255;
    SINE_LUT[424]  = 8'd255;
    SINE_LUT[425]  = 8'd255;
    SINE_LUT[426]  = 8'd255;
    SINE_LUT[427]  = 8'd255;
    SINE_LUT[428]  = 8'd255;
    SINE_LUT[429]  = 8'd255;
    SINE_LUT[430]  = 8'd255;
    SINE_LUT[431]  = 8'd255;
    SINE_LUT[432]  = 8'd255;
    SINE_LUT[433]  = 8'd255;
    SINE_LUT[434]  = 8'd255;
    SINE_LUT[435]  = 8'd255;
    SINE_LUT[436]  = 8'd255;
    SINE_LUT[437]  = 8'd255;
    SINE_LUT[438]  = 8'd255;
    SINE_LUT[439]  = 8'd255;
    SINE_LUT[440]  = 8'd255;
    SINE_LUT[441]  = 8'd255;
    SINE_LUT[442]  = 8'd255;
    SINE_LUT[443]  = 8'd255;
    SINE_LUT[444]  = 8'd255;
    SINE_LUT[445]  = 8'd255;
    SINE_LUT[446]  = 8'd255;
    SINE_LUT[447]  = 8'd255;
    SINE_LUT[448]  = 8'd255;
    SINE_LUT[449]  = 8'd255;
    SINE_LUT[450]  = 8'd255;
    SINE_LUT[451]  = 8'd255;
    SINE_LUT[452]  = 8'd255;
    SINE_LUT[453]  = 8'd255;
    SINE_LUT[454]  = 8'd255;
    SINE_LUT[455]  = 8'd255;
    SINE_LUT[456]  = 8'd255;
    SINE_LUT[457]  = 8'd255;
    SINE_LUT[458]  = 8'd255;
    SINE_LUT[459]  = 8'd255;
    SINE_LUT[460]  = 8'd255;
    SINE_LUT[461]  = 8'd255;
    SINE_LUT[462]  = 8'd255;
    SINE_LUT[463]  = 8'd255;
    SINE_LUT[464]  = 8'd255;
    SINE_LUT[465]  = 8'd254;
    SINE_LUT[466]  = 8'd254;
    SINE_LUT[467]  = 8'd254;
    SINE_LUT[468]  = 8'd254;
    SINE_LUT[469]  = 8'd254;
    SINE_LUT[470]  = 8'd254;
    SINE_LUT[471]  = 8'd254;
    SINE_LUT[472]  = 8'd254;
    SINE_LUT[473]  = 8'd254;
    SINE_LUT[474]  = 8'd254;
    SINE_LUT[475]  = 8'd254;
    SINE_LUT[476]  = 8'd254;
    SINE_LUT[477]  = 8'd254;
    SINE_LUT[478]  = 8'd254;
    SINE_LUT[479]  = 8'd254;
    SINE_LUT[480]  = 8'd254;
    SINE_LUT[481]  = 8'd254;
    SINE_LUT[482]  = 8'd254;
    SINE_LUT[483]  = 8'd253;
    SINE_LUT[484]  = 8'd253;
    SINE_LUT[485]  = 8'd253;
    SINE_LUT[486]  = 8'd253;
    SINE_LUT[487]  = 8'd253;
    SINE_LUT[488]  = 8'd253;
    SINE_LUT[489]  = 8'd253;
    SINE_LUT[490]  = 8'd253;
    SINE_LUT[491]  = 8'd253;
    SINE_LUT[492]  = 8'd253;
    SINE_LUT[493]  = 8'd253;
    SINE_LUT[494]  = 8'd253;
    SINE_LUT[495]  = 8'd252;
    SINE_LUT[496]  = 8'd252;
    SINE_LUT[497]  = 8'd252;
    SINE_LUT[498]  = 8'd252;
    SINE_LUT[499]  = 8'd252;
    SINE_LUT[500]  = 8'd252;
    SINE_LUT[501]  = 8'd252;
    SINE_LUT[502]  = 8'd252;
    SINE_LUT[503]  = 8'd252;
    SINE_LUT[504]  = 8'd252;
    SINE_LUT[505]  = 8'd252;
    SINE_LUT[506]  = 8'd251;
    SINE_LUT[507]  = 8'd251;
    SINE_LUT[508]  = 8'd251;
    SINE_LUT[509]  = 8'd251;
    SINE_LUT[510]  = 8'd251;
    SINE_LUT[511]  = 8'd251;
    SINE_LUT[512]  = 8'd251;
    SINE_LUT[513]  = 8'd251;
    SINE_LUT[514]  = 8'd250;
    SINE_LUT[515]  = 8'd250;
    SINE_LUT[516]  = 8'd250;
    SINE_LUT[517]  = 8'd250;
    SINE_LUT[518]  = 8'd250;
    SINE_LUT[519]  = 8'd250;
    SINE_LUT[520]  = 8'd250;
    SINE_LUT[521]  = 8'd250;
    SINE_LUT[522]  = 8'd249;
    SINE_LUT[523]  = 8'd249;
    SINE_LUT[524]  = 8'd249;
    SINE_LUT[525]  = 8'd249;
    SINE_LUT[526]  = 8'd249;
    SINE_LUT[527]  = 8'd249;
    SINE_LUT[528]  = 8'd249;
    SINE_LUT[529]  = 8'd249;
    SINE_LUT[530]  = 8'd248;
    SINE_LUT[531]  = 8'd248;
    SINE_LUT[532]  = 8'd248;
    SINE_LUT[533]  = 8'd248;
    SINE_LUT[534]  = 8'd248;
    SINE_LUT[535]  = 8'd248;
    SINE_LUT[536]  = 8'd247;
    SINE_LUT[537]  = 8'd247;
    SINE_LUT[538]  = 8'd247;
    SINE_LUT[539]  = 8'd247;
    SINE_LUT[540]  = 8'd247;
    SINE_LUT[541]  = 8'd247;
    SINE_LUT[542]  = 8'd247;
    SINE_LUT[543]  = 8'd246;
    SINE_LUT[544]  = 8'd246;
    SINE_LUT[545]  = 8'd246;
    SINE_LUT[546]  = 8'd246;
    SINE_LUT[547]  = 8'd246;
    SINE_LUT[548]  = 8'd246;
    SINE_LUT[549]  = 8'd245;
    SINE_LUT[550]  = 8'd245;
    SINE_LUT[551]  = 8'd245;
    SINE_LUT[552]  = 8'd245;
    SINE_LUT[553]  = 8'd245;
    SINE_LUT[554]  = 8'd244;
    SINE_LUT[555]  = 8'd244;
    SINE_LUT[556]  = 8'd244;
    SINE_LUT[557]  = 8'd244;
    SINE_LUT[558]  = 8'd244;
    SINE_LUT[559]  = 8'd244;
    SINE_LUT[560]  = 8'd243;
    SINE_LUT[561]  = 8'd243;
    SINE_LUT[562]  = 8'd243;
    SINE_LUT[563]  = 8'd243;
    SINE_LUT[564]  = 8'd243;
    SINE_LUT[565]  = 8'd242;
    SINE_LUT[566]  = 8'd242;
    SINE_LUT[567]  = 8'd242;
    SINE_LUT[568]  = 8'd242;
    SINE_LUT[569]  = 8'd242;
    SINE_LUT[570]  = 8'd241;
    SINE_LUT[571]  = 8'd241;
    SINE_LUT[572]  = 8'd241;
    SINE_LUT[573]  = 8'd241;
    SINE_LUT[574]  = 8'd241;
    SINE_LUT[575]  = 8'd240;
    SINE_LUT[576]  = 8'd240;
    SINE_LUT[577]  = 8'd240;
    SINE_LUT[578]  = 8'd240;
    SINE_LUT[579]  = 8'd239;
    SINE_LUT[580]  = 8'd239;
    SINE_LUT[581]  = 8'd239;
    SINE_LUT[582]  = 8'd239;
    SINE_LUT[583]  = 8'd239;
    SINE_LUT[584]  = 8'd238;
    SINE_LUT[585]  = 8'd238;
    SINE_LUT[586]  = 8'd238;
    SINE_LUT[587]  = 8'd238;
    SINE_LUT[588]  = 8'd237;
    SINE_LUT[589]  = 8'd237;
    SINE_LUT[590]  = 8'd237;
    SINE_LUT[591]  = 8'd237;
    SINE_LUT[592]  = 8'd237;
    SINE_LUT[593]  = 8'd236;
    SINE_LUT[594]  = 8'd236;
    SINE_LUT[595]  = 8'd236;
    SINE_LUT[596]  = 8'd236;
    SINE_LUT[597]  = 8'd235;
    SINE_LUT[598]  = 8'd235;
    SINE_LUT[599]  = 8'd235;
    SINE_LUT[600]  = 8'd235;
    SINE_LUT[601]  = 8'd234;
    SINE_LUT[602]  = 8'd234;
    SINE_LUT[603]  = 8'd234;
    SINE_LUT[604]  = 8'd234;
    SINE_LUT[605]  = 8'd233;
    SINE_LUT[606]  = 8'd233;
    SINE_LUT[607]  = 8'd233;
    SINE_LUT[608]  = 8'd233;
    SINE_LUT[609]  = 8'd232;
    SINE_LUT[610]  = 8'd232;
    SINE_LUT[611]  = 8'd232;
    SINE_LUT[612]  = 8'd232;
    SINE_LUT[613]  = 8'd231;
    SINE_LUT[614]  = 8'd231;
    SINE_LUT[615]  = 8'd231;
    SINE_LUT[616]  = 8'd230;
    SINE_LUT[617]  = 8'd230;
    SINE_LUT[618]  = 8'd230;
    SINE_LUT[619]  = 8'd230;
    SINE_LUT[620]  = 8'd229;
    SINE_LUT[621]  = 8'd229;
    SINE_LUT[622]  = 8'd229;
    SINE_LUT[623]  = 8'd229;
    SINE_LUT[624]  = 8'd228;
    SINE_LUT[625]  = 8'd228;
    SINE_LUT[626]  = 8'd228;
    SINE_LUT[627]  = 8'd227;
    SINE_LUT[628]  = 8'd227;
    SINE_LUT[629]  = 8'd227;
    SINE_LUT[630]  = 8'd227;
    SINE_LUT[631]  = 8'd226;
    SINE_LUT[632]  = 8'd226;
    SINE_LUT[633]  = 8'd226;
    SINE_LUT[634]  = 8'd225;
    SINE_LUT[635]  = 8'd225;
    SINE_LUT[636]  = 8'd225;
    SINE_LUT[637]  = 8'd225;
    SINE_LUT[638]  = 8'd224;
    SINE_LUT[639]  = 8'd224;
    SINE_LUT[640]  = 8'd224;
    SINE_LUT[641]  = 8'd223;
    SINE_LUT[642]  = 8'd223;
    SINE_LUT[643]  = 8'd223;
    SINE_LUT[644]  = 8'd222;
    SINE_LUT[645]  = 8'd222;
    SINE_LUT[646]  = 8'd222;
    SINE_LUT[647]  = 8'd222;
    SINE_LUT[648]  = 8'd221;
    SINE_LUT[649]  = 8'd221;
    SINE_LUT[650]  = 8'd221;
    SINE_LUT[651]  = 8'd220;
    SINE_LUT[652]  = 8'd220;
    SINE_LUT[653]  = 8'd220;
    SINE_LUT[654]  = 8'd219;
    SINE_LUT[655]  = 8'd219;
    SINE_LUT[656]  = 8'd219;
    SINE_LUT[657]  = 8'd218;
    SINE_LUT[658]  = 8'd218;
    SINE_LUT[659]  = 8'd218;
    SINE_LUT[660]  = 8'd217;
    SINE_LUT[661]  = 8'd217;
    SINE_LUT[662]  = 8'd217;
    SINE_LUT[663]  = 8'd216;
    SINE_LUT[664]  = 8'd216;
    SINE_LUT[665]  = 8'd216;
    SINE_LUT[666]  = 8'd215;
    SINE_LUT[667]  = 8'd215;
    SINE_LUT[668]  = 8'd215;
    SINE_LUT[669]  = 8'd214;
    SINE_LUT[670]  = 8'd214;
    SINE_LUT[671]  = 8'd214;
    SINE_LUT[672]  = 8'd213;
    SINE_LUT[673]  = 8'd213;
    SINE_LUT[674]  = 8'd213;
    SINE_LUT[675]  = 8'd212;
    SINE_LUT[676]  = 8'd212;
    SINE_LUT[677]  = 8'd212;
    SINE_LUT[678]  = 8'd211;
    SINE_LUT[679]  = 8'd211;
    SINE_LUT[680]  = 8'd211;
    SINE_LUT[681]  = 8'd210;
    SINE_LUT[682]  = 8'd210;
    SINE_LUT[683]  = 8'd210;
    SINE_LUT[684]  = 8'd209;
    SINE_LUT[685]  = 8'd209;
    SINE_LUT[686]  = 8'd209;
    SINE_LUT[687]  = 8'd208;
    SINE_LUT[688]  = 8'd208;
    SINE_LUT[689]  = 8'd208;
    SINE_LUT[690]  = 8'd207;
    SINE_LUT[691]  = 8'd207;
    SINE_LUT[692]  = 8'd207;
    SINE_LUT[693]  = 8'd206;
    SINE_LUT[694]  = 8'd206;
    SINE_LUT[695]  = 8'd205;
    SINE_LUT[696]  = 8'd205;
    SINE_LUT[697]  = 8'd205;
    SINE_LUT[698]  = 8'd204;
    SINE_LUT[699]  = 8'd204;
    SINE_LUT[700]  = 8'd204;
    SINE_LUT[701]  = 8'd203;
    SINE_LUT[702]  = 8'd203;
    SINE_LUT[703]  = 8'd203;
    SINE_LUT[704]  = 8'd202;
    SINE_LUT[705]  = 8'd202;
    SINE_LUT[706]  = 8'd201;
    SINE_LUT[707]  = 8'd201;
    SINE_LUT[708]  = 8'd201;
    SINE_LUT[709]  = 8'd200;
    SINE_LUT[710]  = 8'd200;
    SINE_LUT[711]  = 8'd200;
    SINE_LUT[712]  = 8'd199;
    SINE_LUT[713]  = 8'd199;
    SINE_LUT[714]  = 8'd198;
    SINE_LUT[715]  = 8'd198;
    SINE_LUT[716]  = 8'd198;
    SINE_LUT[717]  = 8'd197;
    SINE_LUT[718]  = 8'd197;
    SINE_LUT[719]  = 8'd197;
    SINE_LUT[720]  = 8'd196;
    SINE_LUT[721]  = 8'd196;
    SINE_LUT[722]  = 8'd195;
    SINE_LUT[723]  = 8'd195;
    SINE_LUT[724]  = 8'd195;
    SINE_LUT[725]  = 8'd194;
    SINE_LUT[726]  = 8'd194;
    SINE_LUT[727]  = 8'd193;
    SINE_LUT[728]  = 8'd193;
    SINE_LUT[729]  = 8'd193;
    SINE_LUT[730]  = 8'd192;
    SINE_LUT[731]  = 8'd192;
    SINE_LUT[732]  = 8'd192;
    SINE_LUT[733]  = 8'd191;
    SINE_LUT[734]  = 8'd191;
    SINE_LUT[735]  = 8'd190;
    SINE_LUT[736]  = 8'd190;
    SINE_LUT[737]  = 8'd190;
    SINE_LUT[738]  = 8'd189;
    SINE_LUT[739]  = 8'd189;
    SINE_LUT[740]  = 8'd188;
    SINE_LUT[741]  = 8'd188;
    SINE_LUT[742]  = 8'd188;
    SINE_LUT[743]  = 8'd187;
    SINE_LUT[744]  = 8'd187;
    SINE_LUT[745]  = 8'd186;
    SINE_LUT[746]  = 8'd186;
    SINE_LUT[747]  = 8'd186;
    SINE_LUT[748]  = 8'd185;
    SINE_LUT[749]  = 8'd185;
    SINE_LUT[750]  = 8'd184;
    SINE_LUT[751]  = 8'd184;
    SINE_LUT[752]  = 8'd184;
    SINE_LUT[753]  = 8'd183;
    SINE_LUT[754]  = 8'd183;
    SINE_LUT[755]  = 8'd182;
    SINE_LUT[756]  = 8'd182;
    SINE_LUT[757]  = 8'd181;
    SINE_LUT[758]  = 8'd181;
    SINE_LUT[759]  = 8'd181;
    SINE_LUT[760]  = 8'd180;
    SINE_LUT[761]  = 8'd180;
    SINE_LUT[762]  = 8'd179;
    SINE_LUT[763]  = 8'd179;
    SINE_LUT[764]  = 8'd179;
    SINE_LUT[765]  = 8'd178;
    SINE_LUT[766]  = 8'd178;
    SINE_LUT[767]  = 8'd177;
    SINE_LUT[768]  = 8'd177;
    SINE_LUT[769]  = 8'd176;
    SINE_LUT[770]  = 8'd176;
    SINE_LUT[771]  = 8'd176;
    SINE_LUT[772]  = 8'd175;
    SINE_LUT[773]  = 8'd175;
    SINE_LUT[774]  = 8'd174;
    SINE_LUT[775]  = 8'd174;
    SINE_LUT[776]  = 8'd174;
    SINE_LUT[777]  = 8'd173;
    SINE_LUT[778]  = 8'd173;
    SINE_LUT[779]  = 8'd172;
    SINE_LUT[780]  = 8'd172;
    SINE_LUT[781]  = 8'd171;
    SINE_LUT[782]  = 8'd171;
    SINE_LUT[783]  = 8'd171;
    SINE_LUT[784]  = 8'd170;
    SINE_LUT[785]  = 8'd170;
    SINE_LUT[786]  = 8'd169;
    SINE_LUT[787]  = 8'd169;
    SINE_LUT[788]  = 8'd168;
    SINE_LUT[789]  = 8'd168;
    SINE_LUT[790]  = 8'd168;
    SINE_LUT[791]  = 8'd167;
    SINE_LUT[792]  = 8'd167;
    SINE_LUT[793]  = 8'd166;
    SINE_LUT[794]  = 8'd166;
    SINE_LUT[795]  = 8'd165;
    SINE_LUT[796]  = 8'd165;
    SINE_LUT[797]  = 8'd164;
    SINE_LUT[798]  = 8'd164;
    SINE_LUT[799]  = 8'd164;
    SINE_LUT[800]  = 8'd163;
    SINE_LUT[801]  = 8'd163;
    SINE_LUT[802]  = 8'd162;
    SINE_LUT[803]  = 8'd162;
    SINE_LUT[804]  = 8'd161;
    SINE_LUT[805]  = 8'd161;
    SINE_LUT[806]  = 8'd161;
    SINE_LUT[807]  = 8'd160;
    SINE_LUT[808]  = 8'd160;
    SINE_LUT[809]  = 8'd159;
    SINE_LUT[810]  = 8'd159;
    SINE_LUT[811]  = 8'd158;
    SINE_LUT[812]  = 8'd158;
    SINE_LUT[813]  = 8'd157;
    SINE_LUT[814]  = 8'd157;
    SINE_LUT[815]  = 8'd157;
    SINE_LUT[816]  = 8'd156;
    SINE_LUT[817]  = 8'd156;
    SINE_LUT[818]  = 8'd155;
    SINE_LUT[819]  = 8'd155;
    SINE_LUT[820]  = 8'd154;
    SINE_LUT[821]  = 8'd154;
    SINE_LUT[822]  = 8'd153;
    SINE_LUT[823]  = 8'd153;
    SINE_LUT[824]  = 8'd153;
    SINE_LUT[825]  = 8'd152;
    SINE_LUT[826]  = 8'd152;
    SINE_LUT[827]  = 8'd151;
    SINE_LUT[828]  = 8'd151;
    SINE_LUT[829]  = 8'd150;
    SINE_LUT[830]  = 8'd150;
    SINE_LUT[831]  = 8'd149;
    SINE_LUT[832]  = 8'd149;
    SINE_LUT[833]  = 8'd149;
    SINE_LUT[834]  = 8'd148;
    SINE_LUT[835]  = 8'd148;
    SINE_LUT[836]  = 8'd147;
    SINE_LUT[837]  = 8'd147;
    SINE_LUT[838]  = 8'd146;
    SINE_LUT[839]  = 8'd146;
    SINE_LUT[840]  = 8'd145;
    SINE_LUT[841]  = 8'd145;
    SINE_LUT[842]  = 8'd145;
    SINE_LUT[843]  = 8'd144;
    SINE_LUT[844]  = 8'd144;
    SINE_LUT[845]  = 8'd143;
    SINE_LUT[846]  = 8'd143;
    SINE_LUT[847]  = 8'd142;
    SINE_LUT[848]  = 8'd142;
    SINE_LUT[849]  = 8'd141;
    SINE_LUT[850]  = 8'd141;
    SINE_LUT[851]  = 8'd140;
    SINE_LUT[852]  = 8'd140;
    SINE_LUT[853]  = 8'd140;
    SINE_LUT[854]  = 8'd139;
    SINE_LUT[855]  = 8'd139;
    SINE_LUT[856]  = 8'd138;
    SINE_LUT[857]  = 8'd138;
    SINE_LUT[858]  = 8'd137;
    SINE_LUT[859]  = 8'd137;
    SINE_LUT[860]  = 8'd136;
    SINE_LUT[861]  = 8'd136;
    SINE_LUT[862]  = 8'd135;
    SINE_LUT[863]  = 8'd135;
    SINE_LUT[864]  = 8'd135;
    SINE_LUT[865]  = 8'd134;
    SINE_LUT[866]  = 8'd134;
    SINE_LUT[867]  = 8'd133;
    SINE_LUT[868]  = 8'd133;
    SINE_LUT[869]  = 8'd132;
    SINE_LUT[870]  = 8'd132;
    SINE_LUT[871]  = 8'd131;
    SINE_LUT[872]  = 8'd131;
    SINE_LUT[873]  = 8'd130;
    SINE_LUT[874]  = 8'd130;
    SINE_LUT[875]  = 8'd130;
    SINE_LUT[876]  = 8'd129;
    SINE_LUT[877]  = 8'd129;
    SINE_LUT[878]  = 8'd128;
    SINE_LUT[879]  = 8'd128;
    SINE_LUT[880]  = 8'd127;
    SINE_LUT[881]  = 8'd127;
    SINE_LUT[882]  = 8'd126;
    SINE_LUT[883]  = 8'd126;
    SINE_LUT[884]  = 8'd126;
    SINE_LUT[885]  = 8'd125;
    SINE_LUT[886]  = 8'd125;
    SINE_LUT[887]  = 8'd124;
    SINE_LUT[888]  = 8'd124;
    SINE_LUT[889]  = 8'd123;
    SINE_LUT[890]  = 8'd123;
    SINE_LUT[891]  = 8'd122;
    SINE_LUT[892]  = 8'd122;
    SINE_LUT[893]  = 8'd121;
    SINE_LUT[894]  = 8'd121;
    SINE_LUT[895]  = 8'd121;
    SINE_LUT[896]  = 8'd120;
    SINE_LUT[897]  = 8'd120;
    SINE_LUT[898]  = 8'd119;
    SINE_LUT[899]  = 8'd119;
    SINE_LUT[900]  = 8'd118;
    SINE_LUT[901]  = 8'd118;
    SINE_LUT[902]  = 8'd117;
    SINE_LUT[903]  = 8'd117;
    SINE_LUT[904]  = 8'd116;
    SINE_LUT[905]  = 8'd116;
    SINE_LUT[906]  = 8'd116;
    SINE_LUT[907]  = 8'd115;
    SINE_LUT[908]  = 8'd115;
    SINE_LUT[909]  = 8'd114;
    SINE_LUT[910]  = 8'd114;
    SINE_LUT[911]  = 8'd113;
    SINE_LUT[912]  = 8'd113;
    SINE_LUT[913]  = 8'd112;
    SINE_LUT[914]  = 8'd112;
    SINE_LUT[915]  = 8'd111;
    SINE_LUT[916]  = 8'd111;
    SINE_LUT[917]  = 8'd111;
    SINE_LUT[918]  = 8'd110;
    SINE_LUT[919]  = 8'd110;
    SINE_LUT[920]  = 8'd109;
    SINE_LUT[921]  = 8'd109;
    SINE_LUT[922]  = 8'd108;
    SINE_LUT[923]  = 8'd108;
    SINE_LUT[924]  = 8'd107;
    SINE_LUT[925]  = 8'd107;
    SINE_LUT[926]  = 8'd107;
    SINE_LUT[927]  = 8'd106;
    SINE_LUT[928]  = 8'd106;
    SINE_LUT[929]  = 8'd105;
    SINE_LUT[930]  = 8'd105;
    SINE_LUT[931]  = 8'd104;
    SINE_LUT[932]  = 8'd104;
    SINE_LUT[933]  = 8'd103;
    SINE_LUT[934]  = 8'd103;
    SINE_LUT[935]  = 8'd103;
    SINE_LUT[936]  = 8'd102;
    SINE_LUT[937]  = 8'd102;
    SINE_LUT[938]  = 8'd101;
    SINE_LUT[939]  = 8'd101;
    SINE_LUT[940]  = 8'd100;
    SINE_LUT[941]  = 8'd100;
    SINE_LUT[942]  = 8'd99;
    SINE_LUT[943]  = 8'd99;
    SINE_LUT[944]  = 8'd99;
    SINE_LUT[945]  = 8'd98;
    SINE_LUT[946]  = 8'd98;
    SINE_LUT[947]  = 8'd97;
    SINE_LUT[948]  = 8'd97;
    SINE_LUT[949]  = 8'd96;
    SINE_LUT[950]  = 8'd96;
    SINE_LUT[951]  = 8'd95;
    SINE_LUT[952]  = 8'd95;
    SINE_LUT[953]  = 8'd95;
    SINE_LUT[954]  = 8'd94;
    SINE_LUT[955]  = 8'd94;
    SINE_LUT[956]  = 8'd93;
    SINE_LUT[957]  = 8'd93;
    SINE_LUT[958]  = 8'd92;
    SINE_LUT[959]  = 8'd92;
    SINE_LUT[960]  = 8'd92;
    SINE_LUT[961]  = 8'd91;
    SINE_LUT[962]  = 8'd91;
    SINE_LUT[963]  = 8'd90;
    SINE_LUT[964]  = 8'd90;
    SINE_LUT[965]  = 8'd89;
    SINE_LUT[966]  = 8'd89;
    SINE_LUT[967]  = 8'd88;
    SINE_LUT[968]  = 8'd88;
    SINE_LUT[969]  = 8'd88;
    SINE_LUT[970]  = 8'd87;
    SINE_LUT[971]  = 8'd87;
    SINE_LUT[972]  = 8'd86;
    SINE_LUT[973]  = 8'd86;
    SINE_LUT[974]  = 8'd85;
    SINE_LUT[975]  = 8'd85;
    SINE_LUT[976]  = 8'd85;
    SINE_LUT[977]  = 8'd84;
    SINE_LUT[978]  = 8'd84;
    SINE_LUT[979]  = 8'd83;
    SINE_LUT[980]  = 8'd83;
    SINE_LUT[981]  = 8'd82;
    SINE_LUT[982]  = 8'd82;
    SINE_LUT[983]  = 8'd82;
    SINE_LUT[984]  = 8'd81;
    SINE_LUT[985]  = 8'd81;
    SINE_LUT[986]  = 8'd80;
    SINE_LUT[987]  = 8'd80;
    SINE_LUT[988]  = 8'd80;
    SINE_LUT[989]  = 8'd79;
    SINE_LUT[990]  = 8'd79;
    SINE_LUT[991]  = 8'd78;
    SINE_LUT[992]  = 8'd78;
    SINE_LUT[993]  = 8'd77;
    SINE_LUT[994]  = 8'd77;
    SINE_LUT[995]  = 8'd77;
    SINE_LUT[996]  = 8'd76;
    SINE_LUT[997]  = 8'd76;
    SINE_LUT[998]  = 8'd75;
    SINE_LUT[999]  = 8'd75;
    SINE_LUT[1000]  = 8'd75;
    SINE_LUT[1001]  = 8'd74;
    SINE_LUT[1002]  = 8'd74;
    SINE_LUT[1003]  = 8'd73;
    SINE_LUT[1004]  = 8'd73;
    SINE_LUT[1005]  = 8'd72;
    SINE_LUT[1006]  = 8'd72;
    SINE_LUT[1007]  = 8'd72;
    SINE_LUT[1008]  = 8'd71;
    SINE_LUT[1009]  = 8'd71;
    SINE_LUT[1010]  = 8'd70;
    SINE_LUT[1011]  = 8'd70;
    SINE_LUT[1012]  = 8'd70;
    SINE_LUT[1013]  = 8'd69;
    SINE_LUT[1014]  = 8'd69;
    SINE_LUT[1015]  = 8'd68;
    SINE_LUT[1016]  = 8'd68;
    SINE_LUT[1017]  = 8'd68;
    SINE_LUT[1018]  = 8'd67;
    SINE_LUT[1019]  = 8'd67;
    SINE_LUT[1020]  = 8'd66;
    SINE_LUT[1021]  = 8'd66;
    SINE_LUT[1022]  = 8'd66;
    SINE_LUT[1023]  = 8'd65;
    SINE_LUT[1024]  = 8'd65;
    SINE_LUT[1025]  = 8'd64;
    SINE_LUT[1026]  = 8'd64;
    SINE_LUT[1027]  = 8'd64;
    SINE_LUT[1028]  = 8'd63;
    SINE_LUT[1029]  = 8'd63;
    SINE_LUT[1030]  = 8'd63;
    SINE_LUT[1031]  = 8'd62;
    SINE_LUT[1032]  = 8'd62;
    SINE_LUT[1033]  = 8'd61;
    SINE_LUT[1034]  = 8'd61;
    SINE_LUT[1035]  = 8'd61;
    SINE_LUT[1036]  = 8'd60;
    SINE_LUT[1037]  = 8'd60;
    SINE_LUT[1038]  = 8'd59;
    SINE_LUT[1039]  = 8'd59;
    SINE_LUT[1040]  = 8'd59;
    SINE_LUT[1041]  = 8'd58;
    SINE_LUT[1042]  = 8'd58;
    SINE_LUT[1043]  = 8'd58;
    SINE_LUT[1044]  = 8'd57;
    SINE_LUT[1045]  = 8'd57;
    SINE_LUT[1046]  = 8'd56;
    SINE_LUT[1047]  = 8'd56;
    SINE_LUT[1048]  = 8'd56;
    SINE_LUT[1049]  = 8'd55;
    SINE_LUT[1050]  = 8'd55;
    SINE_LUT[1051]  = 8'd55;
    SINE_LUT[1052]  = 8'd54;
    SINE_LUT[1053]  = 8'd54;
    SINE_LUT[1054]  = 8'd53;
    SINE_LUT[1055]  = 8'd53;
    SINE_LUT[1056]  = 8'd53;
    SINE_LUT[1057]  = 8'd52;
    SINE_LUT[1058]  = 8'd52;
    SINE_LUT[1059]  = 8'd52;
    SINE_LUT[1060]  = 8'd51;
    SINE_LUT[1061]  = 8'd51;
    SINE_LUT[1062]  = 8'd51;
    SINE_LUT[1063]  = 8'd50;
    SINE_LUT[1064]  = 8'd50;
    SINE_LUT[1065]  = 8'd49;
    SINE_LUT[1066]  = 8'd49;
    SINE_LUT[1067]  = 8'd49;
    SINE_LUT[1068]  = 8'd48;
    SINE_LUT[1069]  = 8'd48;
    SINE_LUT[1070]  = 8'd48;
    SINE_LUT[1071]  = 8'd47;
    SINE_LUT[1072]  = 8'd47;
    SINE_LUT[1073]  = 8'd47;
    SINE_LUT[1074]  = 8'd46;
    SINE_LUT[1075]  = 8'd46;
    SINE_LUT[1076]  = 8'd46;
    SINE_LUT[1077]  = 8'd45;
    SINE_LUT[1078]  = 8'd45;
    SINE_LUT[1079]  = 8'd45;
    SINE_LUT[1080]  = 8'd44;
    SINE_LUT[1081]  = 8'd44;
    SINE_LUT[1082]  = 8'd44;
    SINE_LUT[1083]  = 8'd43;
    SINE_LUT[1084]  = 8'd43;
    SINE_LUT[1085]  = 8'd43;
    SINE_LUT[1086]  = 8'd42;
    SINE_LUT[1087]  = 8'd42;
    SINE_LUT[1088]  = 8'd42;
    SINE_LUT[1089]  = 8'd41;
    SINE_LUT[1090]  = 8'd41;
    SINE_LUT[1091]  = 8'd41;
    SINE_LUT[1092]  = 8'd40;
    SINE_LUT[1093]  = 8'd40;
    SINE_LUT[1094]  = 8'd40;
    SINE_LUT[1095]  = 8'd39;
    SINE_LUT[1096]  = 8'd39;
    SINE_LUT[1097]  = 8'd39;
    SINE_LUT[1098]  = 8'd38;
    SINE_LUT[1099]  = 8'd38;
    SINE_LUT[1100]  = 8'd38;
    SINE_LUT[1101]  = 8'd37;
    SINE_LUT[1102]  = 8'd37;
    SINE_LUT[1103]  = 8'd37;
    SINE_LUT[1104]  = 8'd36;
    SINE_LUT[1105]  = 8'd36;
    SINE_LUT[1106]  = 8'd36;
    SINE_LUT[1107]  = 8'd35;
    SINE_LUT[1108]  = 8'd35;
    SINE_LUT[1109]  = 8'd35;
    SINE_LUT[1110]  = 8'd34;
    SINE_LUT[1111]  = 8'd34;
    SINE_LUT[1112]  = 8'd34;
    SINE_LUT[1113]  = 8'd34;
    SINE_LUT[1114]  = 8'd33;
    SINE_LUT[1115]  = 8'd33;
    SINE_LUT[1116]  = 8'd33;
    SINE_LUT[1117]  = 8'd32;
    SINE_LUT[1118]  = 8'd32;
    SINE_LUT[1119]  = 8'd32;
    SINE_LUT[1120]  = 8'd31;
    SINE_LUT[1121]  = 8'd31;
    SINE_LUT[1122]  = 8'd31;
    SINE_LUT[1123]  = 8'd31;
    SINE_LUT[1124]  = 8'd30;
    SINE_LUT[1125]  = 8'd30;
    SINE_LUT[1126]  = 8'd30;
    SINE_LUT[1127]  = 8'd29;
    SINE_LUT[1128]  = 8'd29;
    SINE_LUT[1129]  = 8'd29;
    SINE_LUT[1130]  = 8'd29;
    SINE_LUT[1131]  = 8'd28;
    SINE_LUT[1132]  = 8'd28;
    SINE_LUT[1133]  = 8'd28;
    SINE_LUT[1134]  = 8'd27;
    SINE_LUT[1135]  = 8'd27;
    SINE_LUT[1136]  = 8'd27;
    SINE_LUT[1137]  = 8'd27;
    SINE_LUT[1138]  = 8'd26;
    SINE_LUT[1139]  = 8'd26;
    SINE_LUT[1140]  = 8'd26;
    SINE_LUT[1141]  = 8'd26;
    SINE_LUT[1142]  = 8'd25;
    SINE_LUT[1143]  = 8'd25;
    SINE_LUT[1144]  = 8'd25;
    SINE_LUT[1145]  = 8'd24;
    SINE_LUT[1146]  = 8'd24;
    SINE_LUT[1147]  = 8'd24;
    SINE_LUT[1148]  = 8'd24;
    SINE_LUT[1149]  = 8'd23;
    SINE_LUT[1150]  = 8'd23;
    SINE_LUT[1151]  = 8'd23;
    SINE_LUT[1152]  = 8'd23;
    SINE_LUT[1153]  = 8'd22;
    SINE_LUT[1154]  = 8'd22;
    SINE_LUT[1155]  = 8'd22;
    SINE_LUT[1156]  = 8'd22;
    SINE_LUT[1157]  = 8'd21;
    SINE_LUT[1158]  = 8'd21;
    SINE_LUT[1159]  = 8'd21;
    SINE_LUT[1160]  = 8'd21;
    SINE_LUT[1161]  = 8'd20;
    SINE_LUT[1162]  = 8'd20;
    SINE_LUT[1163]  = 8'd20;
    SINE_LUT[1164]  = 8'd20;
    SINE_LUT[1165]  = 8'd19;
    SINE_LUT[1166]  = 8'd19;
    SINE_LUT[1167]  = 8'd19;
    SINE_LUT[1168]  = 8'd19;
    SINE_LUT[1169]  = 8'd19;
    SINE_LUT[1170]  = 8'd18;
    SINE_LUT[1171]  = 8'd18;
    SINE_LUT[1172]  = 8'd18;
    SINE_LUT[1173]  = 8'd18;
    SINE_LUT[1174]  = 8'd17;
    SINE_LUT[1175]  = 8'd17;
    SINE_LUT[1176]  = 8'd17;
    SINE_LUT[1177]  = 8'd17;
    SINE_LUT[1178]  = 8'd17;
    SINE_LUT[1179]  = 8'd16;
    SINE_LUT[1180]  = 8'd16;
    SINE_LUT[1181]  = 8'd16;
    SINE_LUT[1182]  = 8'd16;
    SINE_LUT[1183]  = 8'd15;
    SINE_LUT[1184]  = 8'd15;
    SINE_LUT[1185]  = 8'd15;
    SINE_LUT[1186]  = 8'd15;
    SINE_LUT[1187]  = 8'd15;
    SINE_LUT[1188]  = 8'd14;
    SINE_LUT[1189]  = 8'd14;
    SINE_LUT[1190]  = 8'd14;
    SINE_LUT[1191]  = 8'd14;
    SINE_LUT[1192]  = 8'd14;
    SINE_LUT[1193]  = 8'd13;
    SINE_LUT[1194]  = 8'd13;
    SINE_LUT[1195]  = 8'd13;
    SINE_LUT[1196]  = 8'd13;
    SINE_LUT[1197]  = 8'd13;
    SINE_LUT[1198]  = 8'd12;
    SINE_LUT[1199]  = 8'd12;
    SINE_LUT[1200]  = 8'd12;
    SINE_LUT[1201]  = 8'd12;
    SINE_LUT[1202]  = 8'd12;
    SINE_LUT[1203]  = 8'd12;
    SINE_LUT[1204]  = 8'd11;
    SINE_LUT[1205]  = 8'd11;
    SINE_LUT[1206]  = 8'd11;
    SINE_LUT[1207]  = 8'd11;
    SINE_LUT[1208]  = 8'd11;
    SINE_LUT[1209]  = 8'd10;
    SINE_LUT[1210]  = 8'd10;
    SINE_LUT[1211]  = 8'd10;
    SINE_LUT[1212]  = 8'd10;
    SINE_LUT[1213]  = 8'd10;
    SINE_LUT[1214]  = 8'd10;
    SINE_LUT[1215]  = 8'd9;
    SINE_LUT[1216]  = 8'd9;
    SINE_LUT[1217]  = 8'd9;
    SINE_LUT[1218]  = 8'd9;
    SINE_LUT[1219]  = 8'd9;
    SINE_LUT[1220]  = 8'd9;
    SINE_LUT[1221]  = 8'd9;
    SINE_LUT[1222]  = 8'd8;
    SINE_LUT[1223]  = 8'd8;
    SINE_LUT[1224]  = 8'd8;
    SINE_LUT[1225]  = 8'd8;
    SINE_LUT[1226]  = 8'd8;
    SINE_LUT[1227]  = 8'd8;
    SINE_LUT[1228]  = 8'd7;
    SINE_LUT[1229]  = 8'd7;
    SINE_LUT[1230]  = 8'd7;
    SINE_LUT[1231]  = 8'd7;
    SINE_LUT[1232]  = 8'd7;
    SINE_LUT[1233]  = 8'd7;
    SINE_LUT[1234]  = 8'd7;
    SINE_LUT[1235]  = 8'd7;
    SINE_LUT[1236]  = 8'd6;
    SINE_LUT[1237]  = 8'd6;
    SINE_LUT[1238]  = 8'd6;
    SINE_LUT[1239]  = 8'd6;
    SINE_LUT[1240]  = 8'd6;
    SINE_LUT[1241]  = 8'd6;
    SINE_LUT[1242]  = 8'd6;
    SINE_LUT[1243]  = 8'd6;
    SINE_LUT[1244]  = 8'd5;
    SINE_LUT[1245]  = 8'd5;
    SINE_LUT[1246]  = 8'd5;
    SINE_LUT[1247]  = 8'd5;
    SINE_LUT[1248]  = 8'd5;
    SINE_LUT[1249]  = 8'd5;
    SINE_LUT[1250]  = 8'd5;
    SINE_LUT[1251]  = 8'd5;
    SINE_LUT[1252]  = 8'd4;
    SINE_LUT[1253]  = 8'd4;
    SINE_LUT[1254]  = 8'd4;
    SINE_LUT[1255]  = 8'd4;
    SINE_LUT[1256]  = 8'd4;
    SINE_LUT[1257]  = 8'd4;
    SINE_LUT[1258]  = 8'd4;
    SINE_LUT[1259]  = 8'd4;
    SINE_LUT[1260]  = 8'd4;
    SINE_LUT[1261]  = 8'd4;
    SINE_LUT[1262]  = 8'd4;
    SINE_LUT[1263]  = 8'd3;
    SINE_LUT[1264]  = 8'd3;
    SINE_LUT[1265]  = 8'd3;
    SINE_LUT[1266]  = 8'd3;
    SINE_LUT[1267]  = 8'd3;
    SINE_LUT[1268]  = 8'd3;
    SINE_LUT[1269]  = 8'd3;
    SINE_LUT[1270]  = 8'd3;
    SINE_LUT[1271]  = 8'd3;
    SINE_LUT[1272]  = 8'd3;
    SINE_LUT[1273]  = 8'd3;
    SINE_LUT[1274]  = 8'd3;
    SINE_LUT[1275]  = 8'd2;
    SINE_LUT[1276]  = 8'd2;
    SINE_LUT[1277]  = 8'd2;
    SINE_LUT[1278]  = 8'd2;
    SINE_LUT[1279]  = 8'd2;
    SINE_LUT[1280]  = 8'd2;
    SINE_LUT[1281]  = 8'd2;
    SINE_LUT[1282]  = 8'd2;
    SINE_LUT[1283]  = 8'd2;
    SINE_LUT[1284]  = 8'd2;
    SINE_LUT[1285]  = 8'd2;
    SINE_LUT[1286]  = 8'd2;
    SINE_LUT[1287]  = 8'd2;
    SINE_LUT[1288]  = 8'd2;
    SINE_LUT[1289]  = 8'd2;
    SINE_LUT[1290]  = 8'd2;
    SINE_LUT[1291]  = 8'd2;
    SINE_LUT[1292]  = 8'd2;
    SINE_LUT[1293]  = 8'd1;
    SINE_LUT[1294]  = 8'd1;
    SINE_LUT[1295]  = 8'd1;
    SINE_LUT[1296]  = 8'd1;
    SINE_LUT[1297]  = 8'd1;
    SINE_LUT[1298]  = 8'd1;
    SINE_LUT[1299]  = 8'd1;
    SINE_LUT[1300]  = 8'd1;
    SINE_LUT[1301]  = 8'd1;
    SINE_LUT[1302]  = 8'd1;
    SINE_LUT[1303]  = 8'd1;
    SINE_LUT[1304]  = 8'd1;
    SINE_LUT[1305]  = 8'd1;
    SINE_LUT[1306]  = 8'd1;
    SINE_LUT[1307]  = 8'd1;
    SINE_LUT[1308]  = 8'd1;
    SINE_LUT[1309]  = 8'd1;
    SINE_LUT[1310]  = 8'd1;
    SINE_LUT[1311]  = 8'd1;
    SINE_LUT[1312]  = 8'd1;
    SINE_LUT[1313]  = 8'd1;
    SINE_LUT[1314]  = 8'd1;
    SINE_LUT[1315]  = 8'd1;
    SINE_LUT[1316]  = 8'd1;
    SINE_LUT[1317]  = 8'd1;
    SINE_LUT[1318]  = 8'd1;
    SINE_LUT[1319]  = 8'd1;
    SINE_LUT[1320]  = 8'd1;
    SINE_LUT[1321]  = 8'd1;
    SINE_LUT[1322]  = 8'd1;
    SINE_LUT[1323]  = 8'd1;
    SINE_LUT[1324]  = 8'd1;
    SINE_LUT[1325]  = 8'd1;
    SINE_LUT[1326]  = 8'd1;
    SINE_LUT[1327]  = 8'd1;
    SINE_LUT[1328]  = 8'd1;
    SINE_LUT[1329]  = 8'd1;
    SINE_LUT[1330]  = 8'd1;
    SINE_LUT[1331]  = 8'd1;
    SINE_LUT[1332]  = 8'd1;
    SINE_LUT[1333]  = 8'd1;
    SINE_LUT[1334]  = 8'd1;
    SINE_LUT[1335]  = 8'd1;
    SINE_LUT[1336]  = 8'd1;
    SINE_LUT[1337]  = 8'd1;
    SINE_LUT[1338]  = 8'd1;
    SINE_LUT[1339]  = 8'd1;
    SINE_LUT[1340]  = 8'd1;
    SINE_LUT[1341]  = 8'd1;
    SINE_LUT[1342]  = 8'd1;
    SINE_LUT[1343]  = 8'd2;
    SINE_LUT[1344]  = 8'd2;
    SINE_LUT[1345]  = 8'd2;
    SINE_LUT[1346]  = 8'd2;
    SINE_LUT[1347]  = 8'd2;
    SINE_LUT[1348]  = 8'd2;
    SINE_LUT[1349]  = 8'd2;
    SINE_LUT[1350]  = 8'd2;
    SINE_LUT[1351]  = 8'd2;
    SINE_LUT[1352]  = 8'd2;
    SINE_LUT[1353]  = 8'd2;
    SINE_LUT[1354]  = 8'd2;
    SINE_LUT[1355]  = 8'd2;
    SINE_LUT[1356]  = 8'd2;
    SINE_LUT[1357]  = 8'd2;
    SINE_LUT[1358]  = 8'd2;
    SINE_LUT[1359]  = 8'd2;
    SINE_LUT[1360]  = 8'd2;
    SINE_LUT[1361]  = 8'd3;
    SINE_LUT[1362]  = 8'd3;
    SINE_LUT[1363]  = 8'd3;
    SINE_LUT[1364]  = 8'd3;
    SINE_LUT[1365]  = 8'd3;
    SINE_LUT[1366]  = 8'd3;
    SINE_LUT[1367]  = 8'd3;
    SINE_LUT[1368]  = 8'd3;
    SINE_LUT[1369]  = 8'd3;
    SINE_LUT[1370]  = 8'd3;
    SINE_LUT[1371]  = 8'd3;
    SINE_LUT[1372]  = 8'd3;
    SINE_LUT[1373]  = 8'd3;
    SINE_LUT[1374]  = 8'd4;
    SINE_LUT[1375]  = 8'd4;
    SINE_LUT[1376]  = 8'd4;
    SINE_LUT[1377]  = 8'd4;
    SINE_LUT[1378]  = 8'd4;
    SINE_LUT[1379]  = 8'd4;
    SINE_LUT[1380]  = 8'd4;
    SINE_LUT[1381]  = 8'd4;
    SINE_LUT[1382]  = 8'd4;
    SINE_LUT[1383]  = 8'd4;
    SINE_LUT[1384]  = 8'd5;
    SINE_LUT[1385]  = 8'd5;
    SINE_LUT[1386]  = 8'd5;
    SINE_LUT[1387]  = 8'd5;
    SINE_LUT[1388]  = 8'd5;
    SINE_LUT[1389]  = 8'd5;
    SINE_LUT[1390]  = 8'd5;
    SINE_LUT[1391]  = 8'd5;
    SINE_LUT[1392]  = 8'd5;
    SINE_LUT[1393]  = 8'd6;
    SINE_LUT[1394]  = 8'd6;
    SINE_LUT[1395]  = 8'd6;
    SINE_LUT[1396]  = 8'd6;
    SINE_LUT[1397]  = 8'd6;
    SINE_LUT[1398]  = 8'd6;
    SINE_LUT[1399]  = 8'd6;
    SINE_LUT[1400]  = 8'd6;
    SINE_LUT[1401]  = 8'd7;
    SINE_LUT[1402]  = 8'd7;
    SINE_LUT[1403]  = 8'd7;
    SINE_LUT[1404]  = 8'd7;
    SINE_LUT[1405]  = 8'd7;
    SINE_LUT[1406]  = 8'd7;
    SINE_LUT[1407]  = 8'd7;
    SINE_LUT[1408]  = 8'd8;
    SINE_LUT[1409]  = 8'd8;
    SINE_LUT[1410]  = 8'd8;
    SINE_LUT[1411]  = 8'd8;
    SINE_LUT[1412]  = 8'd8;
    SINE_LUT[1413]  = 8'd8;
    SINE_LUT[1414]  = 8'd8;
    SINE_LUT[1415]  = 8'd9;
    SINE_LUT[1416]  = 8'd9;
    SINE_LUT[1417]  = 8'd9;
    SINE_LUT[1418]  = 8'd9;
    SINE_LUT[1419]  = 8'd9;
    SINE_LUT[1420]  = 8'd9;
    SINE_LUT[1421]  = 8'd10;
    SINE_LUT[1422]  = 8'd10;
    SINE_LUT[1423]  = 8'd10;
    SINE_LUT[1424]  = 8'd10;
    SINE_LUT[1425]  = 8'd10;
    SINE_LUT[1426]  = 8'd10;
    SINE_LUT[1427]  = 8'd11;
    SINE_LUT[1428]  = 8'd11;
    SINE_LUT[1429]  = 8'd11;
    SINE_LUT[1430]  = 8'd11;
    SINE_LUT[1431]  = 8'd11;
    SINE_LUT[1432]  = 8'd11;
    SINE_LUT[1433]  = 8'd12;
    SINE_LUT[1434]  = 8'd12;
    SINE_LUT[1435]  = 8'd12;
    SINE_LUT[1436]  = 8'd12;
    SINE_LUT[1437]  = 8'd12;
    SINE_LUT[1438]  = 8'd13;
    SINE_LUT[1439]  = 8'd13;
    SINE_LUT[1440]  = 8'd13;
    SINE_LUT[1441]  = 8'd13;
    SINE_LUT[1442]  = 8'd13;
    SINE_LUT[1443]  = 8'd14;
    SINE_LUT[1444]  = 8'd14;
    SINE_LUT[1445]  = 8'd14;
    SINE_LUT[1446]  = 8'd14;
    SINE_LUT[1447]  = 8'd14;
    SINE_LUT[1448]  = 8'd15;
    SINE_LUT[1449]  = 8'd15;
    SINE_LUT[1450]  = 8'd15;
    SINE_LUT[1451]  = 8'd15;
    SINE_LUT[1452]  = 8'd15;
    SINE_LUT[1453]  = 8'd16;
    SINE_LUT[1454]  = 8'd16;
    SINE_LUT[1455]  = 8'd16;
    SINE_LUT[1456]  = 8'd16;
    SINE_LUT[1457]  = 8'd16;
    SINE_LUT[1458]  = 8'd17;
    SINE_LUT[1459]  = 8'd17;
    SINE_LUT[1460]  = 8'd17;
    SINE_LUT[1461]  = 8'd17;
    SINE_LUT[1462]  = 8'd18;
    SINE_LUT[1463]  = 8'd18;
    SINE_LUT[1464]  = 8'd18;
    SINE_LUT[1465]  = 8'd18;
    SINE_LUT[1466]  = 8'd18;
    SINE_LUT[1467]  = 8'd19;
    SINE_LUT[1468]  = 8'd19;
    SINE_LUT[1469]  = 8'd19;
    SINE_LUT[1470]  = 8'd19;
    SINE_LUT[1471]  = 8'd20;
    SINE_LUT[1472]  = 8'd20;
    SINE_LUT[1473]  = 8'd20;
    SINE_LUT[1474]  = 8'd20;
    SINE_LUT[1475]  = 8'd21;
    SINE_LUT[1476]  = 8'd21;
    SINE_LUT[1477]  = 8'd21;
    SINE_LUT[1478]  = 8'd21;
    SINE_LUT[1479]  = 8'd22;
    SINE_LUT[1480]  = 8'd22;
    SINE_LUT[1481]  = 8'd22;
    SINE_LUT[1482]  = 8'd22;
    SINE_LUT[1483]  = 8'd23;
    SINE_LUT[1484]  = 8'd23;
    SINE_LUT[1485]  = 8'd23;
    SINE_LUT[1486]  = 8'd23;
    SINE_LUT[1487]  = 8'd24;
    SINE_LUT[1488]  = 8'd24;
    SINE_LUT[1489]  = 8'd24;
    SINE_LUT[1490]  = 8'd24;
    SINE_LUT[1491]  = 8'd25;
    SINE_LUT[1492]  = 8'd25;
    SINE_LUT[1493]  = 8'd25;
    SINE_LUT[1494]  = 8'd25;
    SINE_LUT[1495]  = 8'd26;
    SINE_LUT[1496]  = 8'd26;
    SINE_LUT[1497]  = 8'd26;
    SINE_LUT[1498]  = 8'd26;
    SINE_LUT[1499]  = 8'd27;
    SINE_LUT[1500]  = 8'd27;
    SINE_LUT[1501]  = 8'd27;
    SINE_LUT[1502]  = 8'd28;
    SINE_LUT[1503]  = 8'd28;
    SINE_LUT[1504]  = 8'd28;
    SINE_LUT[1505]  = 8'd28;
    SINE_LUT[1506]  = 8'd29;
    SINE_LUT[1507]  = 8'd29;
    SINE_LUT[1508]  = 8'd29;
    SINE_LUT[1509]  = 8'd30;
    SINE_LUT[1510]  = 8'd30;
    SINE_LUT[1511]  = 8'd30;
    SINE_LUT[1512]  = 8'd30;
    SINE_LUT[1513]  = 8'd31;
    SINE_LUT[1514]  = 8'd31;
    SINE_LUT[1515]  = 8'd31;
    SINE_LUT[1516]  = 8'd32;
    SINE_LUT[1517]  = 8'd32;
    SINE_LUT[1518]  = 8'd32;
    SINE_LUT[1519]  = 8'd32;
    SINE_LUT[1520]  = 8'd33;
    SINE_LUT[1521]  = 8'd33;
    SINE_LUT[1522]  = 8'd33;
    SINE_LUT[1523]  = 8'd34;
    SINE_LUT[1524]  = 8'd34;
    SINE_LUT[1525]  = 8'd34;
    SINE_LUT[1526]  = 8'd35;
    SINE_LUT[1527]  = 8'd35;
    SINE_LUT[1528]  = 8'd35;
    SINE_LUT[1529]  = 8'd36;
    SINE_LUT[1530]  = 8'd36;
    SINE_LUT[1531]  = 8'd36;
    SINE_LUT[1532]  = 8'd36;
    SINE_LUT[1533]  = 8'd37;
    SINE_LUT[1534]  = 8'd37;
    SINE_LUT[1535]  = 8'd37;
    SINE_LUT[1536]  = 8'd38;
    SINE_LUT[1537]  = 8'd38;
    SINE_LUT[1538]  = 8'd38;
    SINE_LUT[1539]  = 8'd39;
    SINE_LUT[1540]  = 8'd39;
    SINE_LUT[1541]  = 8'd39;
    SINE_LUT[1542]  = 8'd40;
    SINE_LUT[1543]  = 8'd40;
    SINE_LUT[1544]  = 8'd40;
    SINE_LUT[1545]  = 8'd41;
    SINE_LUT[1546]  = 8'd41;
    SINE_LUT[1547]  = 8'd41;
    SINE_LUT[1548]  = 8'd42;
    SINE_LUT[1549]  = 8'd42;
    SINE_LUT[1550]  = 8'd42;
    SINE_LUT[1551]  = 8'd43;
    SINE_LUT[1552]  = 8'd43;
    SINE_LUT[1553]  = 8'd43;
    SINE_LUT[1554]  = 8'd44;
    SINE_LUT[1555]  = 8'd44;
    SINE_LUT[1556]  = 8'd44;
    SINE_LUT[1557]  = 8'd45;
    SINE_LUT[1558]  = 8'd45;
    SINE_LUT[1559]  = 8'd45;
    SINE_LUT[1560]  = 8'd46;
    SINE_LUT[1561]  = 8'd46;
    SINE_LUT[1562]  = 8'd46;
    SINE_LUT[1563]  = 8'd47;
    SINE_LUT[1564]  = 8'd47;
    SINE_LUT[1565]  = 8'd47;
    SINE_LUT[1566]  = 8'd48;
    SINE_LUT[1567]  = 8'd48;
    SINE_LUT[1568]  = 8'd49;
    SINE_LUT[1569]  = 8'd49;
    SINE_LUT[1570]  = 8'd49;
    SINE_LUT[1571]  = 8'd50;
    SINE_LUT[1572]  = 8'd50;
    SINE_LUT[1573]  = 8'd50;
    SINE_LUT[1574]  = 8'd51;
    SINE_LUT[1575]  = 8'd51;
    SINE_LUT[1576]  = 8'd51;
    SINE_LUT[1577]  = 8'd52;
    SINE_LUT[1578]  = 8'd52;
    SINE_LUT[1579]  = 8'd53;
    SINE_LUT[1580]  = 8'd53;
    SINE_LUT[1581]  = 8'd53;
    SINE_LUT[1582]  = 8'd54;
    SINE_LUT[1583]  = 8'd54;
    SINE_LUT[1584]  = 8'd54;
    SINE_LUT[1585]  = 8'd55;
    SINE_LUT[1586]  = 8'd55;
    SINE_LUT[1587]  = 8'd55;
    SINE_LUT[1588]  = 8'd56;
    SINE_LUT[1589]  = 8'd56;
    SINE_LUT[1590]  = 8'd57;
    SINE_LUT[1591]  = 8'd57;
    SINE_LUT[1592]  = 8'd57;
    SINE_LUT[1593]  = 8'd58;
    SINE_LUT[1594]  = 8'd58;
    SINE_LUT[1595]  = 8'd58;
    SINE_LUT[1596]  = 8'd59;
    SINE_LUT[1597]  = 8'd59;
    SINE_LUT[1598]  = 8'd60;
    SINE_LUT[1599]  = 8'd60;
    SINE_LUT[1600]  = 8'd60;
    SINE_LUT[1601]  = 8'd61;
    SINE_LUT[1602]  = 8'd61;
    SINE_LUT[1603]  = 8'd62;
    SINE_LUT[1604]  = 8'd62;
    SINE_LUT[1605]  = 8'd62;
    SINE_LUT[1606]  = 8'd63;
    SINE_LUT[1607]  = 8'd63;
    SINE_LUT[1608]  = 8'd63;
    SINE_LUT[1609]  = 8'd64;
    SINE_LUT[1610]  = 8'd64;
    SINE_LUT[1611]  = 8'd65;
    SINE_LUT[1612]  = 8'd65;
    SINE_LUT[1613]  = 8'd65;
    SINE_LUT[1614]  = 8'd66;
    SINE_LUT[1615]  = 8'd66;
    SINE_LUT[1616]  = 8'd67;
    SINE_LUT[1617]  = 8'd67;
    SINE_LUT[1618]  = 8'd67;
    SINE_LUT[1619]  = 8'd68;
    SINE_LUT[1620]  = 8'd68;
    SINE_LUT[1621]  = 8'd69;
    SINE_LUT[1622]  = 8'd69;
    SINE_LUT[1623]  = 8'd69;
    SINE_LUT[1624]  = 8'd70;
    SINE_LUT[1625]  = 8'd70;
    SINE_LUT[1626]  = 8'd71;
    SINE_LUT[1627]  = 8'd71;
    SINE_LUT[1628]  = 8'd71;
    SINE_LUT[1629]  = 8'd72;
    SINE_LUT[1630]  = 8'd72;
    SINE_LUT[1631]  = 8'd73;
    SINE_LUT[1632]  = 8'd73;
    SINE_LUT[1633]  = 8'd74;
    SINE_LUT[1634]  = 8'd74;
    SINE_LUT[1635]  = 8'd74;
    SINE_LUT[1636]  = 8'd75;
    SINE_LUT[1637]  = 8'd75;
    SINE_LUT[1638]  = 8'd76;
    SINE_LUT[1639]  = 8'd76;
    SINE_LUT[1640]  = 8'd76;
    SINE_LUT[1641]  = 8'd77;
    SINE_LUT[1642]  = 8'd77;
    SINE_LUT[1643]  = 8'd78;
    SINE_LUT[1644]  = 8'd78;
    SINE_LUT[1645]  = 8'd78;
    SINE_LUT[1646]  = 8'd79;
    SINE_LUT[1647]  = 8'd79;
    SINE_LUT[1648]  = 8'd80;
    SINE_LUT[1649]  = 8'd80;
    SINE_LUT[1650]  = 8'd81;
    SINE_LUT[1651]  = 8'd81;
    SINE_LUT[1652]  = 8'd81;
    SINE_LUT[1653]  = 8'd82;
    SINE_LUT[1654]  = 8'd82;
    SINE_LUT[1655]  = 8'd83;
    SINE_LUT[1656]  = 8'd83;
    SINE_LUT[1657]  = 8'd84;
    SINE_LUT[1658]  = 8'd84;
    SINE_LUT[1659]  = 8'd84;
    SINE_LUT[1660]  = 8'd85;
    SINE_LUT[1661]  = 8'd85;
    SINE_LUT[1662]  = 8'd86;
    SINE_LUT[1663]  = 8'd86;
    SINE_LUT[1664]  = 8'd87;
    SINE_LUT[1665]  = 8'd87;
    SINE_LUT[1666]  = 8'd87;
    SINE_LUT[1667]  = 8'd88;
    SINE_LUT[1668]  = 8'd88;
    SINE_LUT[1669]  = 8'd89;
    SINE_LUT[1670]  = 8'd89;
    SINE_LUT[1671]  = 8'd90;
    SINE_LUT[1672]  = 8'd90;
    SINE_LUT[1673]  = 8'd90;
    SINE_LUT[1674]  = 8'd91;
    SINE_LUT[1675]  = 8'd91;
    SINE_LUT[1676]  = 8'd92;
    SINE_LUT[1677]  = 8'd92;
    SINE_LUT[1678]  = 8'd93;
    SINE_LUT[1679]  = 8'd93;
    SINE_LUT[1680]  = 8'd93;
    SINE_LUT[1681]  = 8'd94;
    SINE_LUT[1682]  = 8'd94;
    SINE_LUT[1683]  = 8'd95;
    SINE_LUT[1684]  = 8'd95;
    SINE_LUT[1685]  = 8'd96;
    SINE_LUT[1686]  = 8'd96;
    SINE_LUT[1687]  = 8'd97;
    SINE_LUT[1688]  = 8'd97;
    SINE_LUT[1689]  = 8'd97;
    SINE_LUT[1690]  = 8'd98;
    SINE_LUT[1691]  = 8'd98;
    SINE_LUT[1692]  = 8'd99;
    SINE_LUT[1693]  = 8'd99;
    SINE_LUT[1694]  = 8'd100;
    SINE_LUT[1695]  = 8'd100;
    SINE_LUT[1696]  = 8'd101;
    SINE_LUT[1697]  = 8'd101;
    SINE_LUT[1698]  = 8'd101;
    SINE_LUT[1699]  = 8'd102;
    SINE_LUT[1700]  = 8'd102;
    SINE_LUT[1701]  = 8'd103;
    SINE_LUT[1702]  = 8'd103;
    SINE_LUT[1703]  = 8'd104;
    SINE_LUT[1704]  = 8'd104;
    SINE_LUT[1705]  = 8'd105;
    SINE_LUT[1706]  = 8'd105;
    SINE_LUT[1707]  = 8'd105;
    SINE_LUT[1708]  = 8'd106;
    SINE_LUT[1709]  = 8'd106;
    SINE_LUT[1710]  = 8'd107;
    SINE_LUT[1711]  = 8'd107;
    SINE_LUT[1712]  = 8'd108;
    SINE_LUT[1713]  = 8'd108;
    SINE_LUT[1714]  = 8'd109;
    SINE_LUT[1715]  = 8'd109;
    SINE_LUT[1716]  = 8'd109;
    SINE_LUT[1717]  = 8'd110;
    SINE_LUT[1718]  = 8'd110;
    SINE_LUT[1719]  = 8'd111;
    SINE_LUT[1720]  = 8'd111;
    SINE_LUT[1721]  = 8'd112;
    SINE_LUT[1722]  = 8'd112;
    SINE_LUT[1723]  = 8'd113;
    SINE_LUT[1724]  = 8'd113;
    SINE_LUT[1725]  = 8'd113;
    SINE_LUT[1726]  = 8'd114;
    SINE_LUT[1727]  = 8'd114;
    SINE_LUT[1728]  = 8'd115;
    SINE_LUT[1729]  = 8'd115;
    SINE_LUT[1730]  = 8'd116;
    SINE_LUT[1731]  = 8'd116;
    SINE_LUT[1732]  = 8'd117;
    SINE_LUT[1733]  = 8'd117;
    SINE_LUT[1734]  = 8'd118;
    SINE_LUT[1735]  = 8'd118;
    SINE_LUT[1736]  = 8'd118;
    SINE_LUT[1737]  = 8'd119;
    SINE_LUT[1738]  = 8'd119;
    SINE_LUT[1739]  = 8'd120;
    SINE_LUT[1740]  = 8'd120;
    SINE_LUT[1741]  = 8'd121;
    SINE_LUT[1742]  = 8'd121;
    SINE_LUT[1743]  = 8'd122;
    SINE_LUT[1744]  = 8'd122;
    SINE_LUT[1745]  = 8'd123;
    SINE_LUT[1746]  = 8'd123;
    SINE_LUT[1747]  = 8'd123;
    SINE_LUT[1748]  = 8'd124;
    SINE_LUT[1749]  = 8'd124;
    SINE_LUT[1750]  = 8'd125;
    SINE_LUT[1751]  = 8'd125;
    SINE_LUT[1752]  = 8'd126;
    SINE_LUT[1753]  = 8'd126;
    SINE_LUT[1754]  = 8'd127;
    SINE_LUT[1755]  = 8'd127;
    SINE_LUT[1756]  = 8'd128;
end

  //——— phase pointer & wrap-around logic ———————————
  logic [11:0] ptr;
  logic [11:0] nxt;

  always_ff @(posedge clk or posedge rst) begin
    if (rst)
      ptr <= '0;
    else if (in_valid) begin
      // compute next pointer, with wrap at MAX_INDEX+1
      nxt = ptr + STEP_LUT[in_data];
      if (nxt > 1756)
        ptr <= nxt - (1756 + 1);
      else
        ptr <= nxt;
    end
  end

  //——— output from sine table ————————————————
  assign out_data = SINE_LUT[ptr];
  
endmodule
