module triangle_wave_gen_d (
    input  logic        clk,       // your 50 MHz clock
    input  logic        rst,     
    input  logic        in_valid,  // pulse when new rx_data sample is ready
    input  logic [7:0]  in_data,       // 0–255 sine input
    output logic [7:0]  out_data
);

    // ----------------------------------------------------------------
    // Triangle Lookup Table (user-generated)
    // ----------------------------------------------------------------
    logic [7:0] TRI_LUT [0:500];
    logic [8:0] ptr;
    logic [8:0] nxt;

initial begin
    TRI_LUT[0]  = 8'd128;
    TRI_LUT[1]  = 8'd129;
    TRI_LUT[2]  = 8'd130;
    TRI_LUT[3]  = 8'd131;
    TRI_LUT[4]  = 8'd132;
    TRI_LUT[5]  = 8'd133;
    TRI_LUT[6]  = 8'd134;
    TRI_LUT[7]  = 8'd135;
    TRI_LUT[8]  = 8'd136;
    TRI_LUT[9]  = 8'd137;
    TRI_LUT[10]  = 8'd138;
    TRI_LUT[11]  = 8'd139;
    TRI_LUT[12]  = 8'd140;
    TRI_LUT[13]  = 8'd141;
    TRI_LUT[14]  = 8'd142;
    TRI_LUT[15]  = 8'd143;
    TRI_LUT[16]  = 8'd144;
    TRI_LUT[17]  = 8'd145;
    TRI_LUT[18]  = 8'd146;
    TRI_LUT[19]  = 8'd147;
    TRI_LUT[20]  = 8'd148;
    TRI_LUT[21]  = 8'd149;
    TRI_LUT[22]  = 8'd150;
    TRI_LUT[23]  = 8'd151;
    TRI_LUT[24]  = 8'd152;
    TRI_LUT[25]  = 8'd153;
    TRI_LUT[26]  = 8'd154;
    TRI_LUT[27]  = 8'd155;
    TRI_LUT[28]  = 8'd156;
    TRI_LUT[29]  = 8'd157;
    TRI_LUT[30]  = 8'd158;
    TRI_LUT[31]  = 8'd159;
    TRI_LUT[32]  = 8'd160;
    TRI_LUT[33]  = 8'd161;
    TRI_LUT[34]  = 8'd162;
    TRI_LUT[35]  = 8'd163;
    TRI_LUT[36]  = 8'd165;
    TRI_LUT[37]  = 8'd166;
    TRI_LUT[38]  = 8'd167;
    TRI_LUT[39]  = 8'd168;
    TRI_LUT[40]  = 8'd169;
    TRI_LUT[41]  = 8'd170;
    TRI_LUT[42]  = 8'd171;
    TRI_LUT[43]  = 8'd172;
    TRI_LUT[44]  = 8'd173;
    TRI_LUT[45]  = 8'd174;
    TRI_LUT[46]  = 8'd175;
    TRI_LUT[47]  = 8'd176;
    TRI_LUT[48]  = 8'd177;
    TRI_LUT[49]  = 8'd178;
    TRI_LUT[50]  = 8'd179;
    TRI_LUT[51]  = 8'd180;
    TRI_LUT[52]  = 8'd181;
    TRI_LUT[53]  = 8'd182;
    TRI_LUT[54]  = 8'd183;
    TRI_LUT[55]  = 8'd184;
    TRI_LUT[56]  = 8'd185;
    TRI_LUT[57]  = 8'd186;
    TRI_LUT[58]  = 8'd187;
    TRI_LUT[59]  = 8'd188;
    TRI_LUT[60]  = 8'd189;
    TRI_LUT[61]  = 8'd190;
    TRI_LUT[62]  = 8'd191;
    TRI_LUT[63]  = 8'd192;
    TRI_LUT[64]  = 8'd193;
    TRI_LUT[65]  = 8'd194;
    TRI_LUT[66]  = 8'd195;
    TRI_LUT[67]  = 8'd196;
    TRI_LUT[68]  = 8'd197;
    TRI_LUT[69]  = 8'd198;
    TRI_LUT[70]  = 8'd199;
    TRI_LUT[71]  = 8'd200;
    TRI_LUT[72]  = 8'd201;
    TRI_LUT[73]  = 8'd202;
    TRI_LUT[74]  = 8'd203;
    TRI_LUT[75]  = 8'd204;
    TRI_LUT[76]  = 8'd205;
    TRI_LUT[77]  = 8'd206;
    TRI_LUT[78]  = 8'd207;
    TRI_LUT[79]  = 8'd208;
    TRI_LUT[80]  = 8'd209;
    TRI_LUT[81]  = 8'd210;
    TRI_LUT[82]  = 8'd211;
    TRI_LUT[83]  = 8'd212;
    TRI_LUT[84]  = 8'd213;
    TRI_LUT[85]  = 8'd214;
    TRI_LUT[86]  = 8'd215;
    TRI_LUT[87]  = 8'd216;
    TRI_LUT[88]  = 8'd217;
    TRI_LUT[89]  = 8'd218;
    TRI_LUT[90]  = 8'd219;
    TRI_LUT[91]  = 8'd220;
    TRI_LUT[92]  = 8'd221;
    TRI_LUT[93]  = 8'd222;
    TRI_LUT[94]  = 8'd223;
    TRI_LUT[95]  = 8'd224;
    TRI_LUT[96]  = 8'd225;
    TRI_LUT[97]  = 8'd226;
    TRI_LUT[98]  = 8'd227;
    TRI_LUT[99]  = 8'd228;
    TRI_LUT[100]  = 8'd229;
    TRI_LUT[101]  = 8'd230;
    TRI_LUT[102]  = 8'd231;
    TRI_LUT[103]  = 8'd232;
    TRI_LUT[104]  = 8'd233;
    TRI_LUT[105]  = 8'd234;
    TRI_LUT[106]  = 8'd235;
    TRI_LUT[107]  = 8'd236;
    TRI_LUT[108]  = 8'd238;
    TRI_LUT[109]  = 8'd239;
    TRI_LUT[110]  = 8'd240;
    TRI_LUT[111]  = 8'd241;
    TRI_LUT[112]  = 8'd242;
    TRI_LUT[113]  = 8'd243;
    TRI_LUT[114]  = 8'd244;
    TRI_LUT[115]  = 8'd245;
    TRI_LUT[116]  = 8'd246;
    TRI_LUT[117]  = 8'd247;
    TRI_LUT[118]  = 8'd248;
    TRI_LUT[119]  = 8'd249;
    TRI_LUT[120]  = 8'd250;
    TRI_LUT[121]  = 8'd251;
    TRI_LUT[122]  = 8'd252;
    TRI_LUT[123]  = 8'd253;
    TRI_LUT[124]  = 8'd254;
    TRI_LUT[125]  = 8'd255;
    TRI_LUT[126]  = 8'd254;
    TRI_LUT[127]  = 8'd253;
    TRI_LUT[128]  = 8'd252;
    TRI_LUT[129]  = 8'd251;
    TRI_LUT[130]  = 8'd250;
    TRI_LUT[131]  = 8'd249;
    TRI_LUT[132]  = 8'd248;
    TRI_LUT[133]  = 8'd247;
    TRI_LUT[134]  = 8'd246;
    TRI_LUT[135]  = 8'd245;
    TRI_LUT[136]  = 8'd244;
    TRI_LUT[137]  = 8'd243;
    TRI_LUT[138]  = 8'd242;
    TRI_LUT[139]  = 8'd241;
    TRI_LUT[140]  = 8'd240;
    TRI_LUT[141]  = 8'd239;
    TRI_LUT[142]  = 8'd238;
    TRI_LUT[143]  = 8'd237;
    TRI_LUT[144]  = 8'd236;
    TRI_LUT[145]  = 8'd235;
    TRI_LUT[146]  = 8'd234;
    TRI_LUT[147]  = 8'd233;
    TRI_LUT[148]  = 8'd232;
    TRI_LUT[149]  = 8'd231;
    TRI_LUT[150]  = 8'd230;
    TRI_LUT[151]  = 8'd229;
    TRI_LUT[152]  = 8'd228;
    TRI_LUT[153]  = 8'd227;
    TRI_LUT[154]  = 8'd226;
    TRI_LUT[155]  = 8'd225;
    TRI_LUT[156]  = 8'd224;
    TRI_LUT[157]  = 8'd223;
    TRI_LUT[158]  = 8'd222;
    TRI_LUT[159]  = 8'd221;
    TRI_LUT[160]  = 8'd220;
    TRI_LUT[161]  = 8'd219;
    TRI_LUT[162]  = 8'd218;
    TRI_LUT[163]  = 8'd217;
    TRI_LUT[164]  = 8'd216;
    TRI_LUT[165]  = 8'd215;
    TRI_LUT[166]  = 8'd214;
    TRI_LUT[167]  = 8'd213;
    TRI_LUT[168]  = 8'd212;
    TRI_LUT[169]  = 8'd211;
    TRI_LUT[170]  = 8'd210;
    TRI_LUT[171]  = 8'd209;
    TRI_LUT[172]  = 8'd208;
    TRI_LUT[173]  = 8'd207;
    TRI_LUT[174]  = 8'd206;
    TRI_LUT[175]  = 8'd205;
    TRI_LUT[176]  = 8'd204;
    TRI_LUT[177]  = 8'd203;
    TRI_LUT[178]  = 8'd202;
    TRI_LUT[179]  = 8'd200;
    TRI_LUT[180]  = 8'd199;
    TRI_LUT[181]  = 8'd198;
    TRI_LUT[182]  = 8'd197;
    TRI_LUT[183]  = 8'd196;
    TRI_LUT[184]  = 8'd195;
    TRI_LUT[185]  = 8'd194;
    TRI_LUT[186]  = 8'd193;
    TRI_LUT[187]  = 8'd192;
    TRI_LUT[188]  = 8'd191;
    TRI_LUT[189]  = 8'd190;
    TRI_LUT[190]  = 8'd189;
    TRI_LUT[191]  = 8'd188;
    TRI_LUT[192]  = 8'd187;
    TRI_LUT[193]  = 8'd186;
    TRI_LUT[194]  = 8'd185;
    TRI_LUT[195]  = 8'd184;
    TRI_LUT[196]  = 8'd183;
    TRI_LUT[197]  = 8'd182;
    TRI_LUT[198]  = 8'd181;
    TRI_LUT[199]  = 8'd180;
    TRI_LUT[200]  = 8'd179;
    TRI_LUT[201]  = 8'd178;
    TRI_LUT[202]  = 8'd177;
    TRI_LUT[203]  = 8'd176;
    TRI_LUT[204]  = 8'd175;
    TRI_LUT[205]  = 8'd174;
    TRI_LUT[206]  = 8'd173;
    TRI_LUT[207]  = 8'd172;
    TRI_LUT[208]  = 8'd171;
    TRI_LUT[209]  = 8'd170;
    TRI_LUT[210]  = 8'd169;
    TRI_LUT[211]  = 8'd168;
    TRI_LUT[212]  = 8'd167;
    TRI_LUT[213]  = 8'd166;
    TRI_LUT[214]  = 8'd165;
    TRI_LUT[215]  = 8'd164;
    TRI_LUT[216]  = 8'd163;
    TRI_LUT[217]  = 8'd162;
    TRI_LUT[218]  = 8'd161;
    TRI_LUT[219]  = 8'd160;
    TRI_LUT[220]  = 8'd159;
    TRI_LUT[221]  = 8'd158;
    TRI_LUT[222]  = 8'd157;
    TRI_LUT[223]  = 8'd156;
    TRI_LUT[224]  = 8'd155;
    TRI_LUT[225]  = 8'd154;
    TRI_LUT[226]  = 8'd153;
    TRI_LUT[227]  = 8'd152;
    TRI_LUT[228]  = 8'd151;
    TRI_LUT[229]  = 8'd150;
    TRI_LUT[230]  = 8'd149;
    TRI_LUT[231]  = 8'd148;
    TRI_LUT[232]  = 8'd147;
    TRI_LUT[233]  = 8'd146;
    TRI_LUT[234]  = 8'd145;
    TRI_LUT[235]  = 8'd144;
    TRI_LUT[236]  = 8'd143;
    TRI_LUT[237]  = 8'd142;
    TRI_LUT[238]  = 8'd141;
    TRI_LUT[239]  = 8'd140;
    TRI_LUT[240]  = 8'd139;
    TRI_LUT[241]  = 8'd138;
    TRI_LUT[242]  = 8'd137;
    TRI_LUT[243]  = 8'd136;
    TRI_LUT[244]  = 8'd135;
    TRI_LUT[245]  = 8'd134;
    TRI_LUT[246]  = 8'd133;
    TRI_LUT[247]  = 8'd132;
    TRI_LUT[248]  = 8'd131;
    TRI_LUT[249]  = 8'd130;
    TRI_LUT[250]  = 8'd129;
    TRI_LUT[251]  = 8'd127;
    TRI_LUT[252]  = 8'd126;
    TRI_LUT[253]  = 8'd125;
    TRI_LUT[254]  = 8'd124;
    TRI_LUT[255]  = 8'd123;
    TRI_LUT[256]  = 8'd122;
    TRI_LUT[257]  = 8'd121;
    TRI_LUT[258]  = 8'd120;
    TRI_LUT[259]  = 8'd119;
    TRI_LUT[260]  = 8'd118;
    TRI_LUT[261]  = 8'd117;
    TRI_LUT[262]  = 8'd116;
    TRI_LUT[263]  = 8'd115;
    TRI_LUT[264]  = 8'd114;
    TRI_LUT[265]  = 8'd113;
    TRI_LUT[266]  = 8'd112;
    TRI_LUT[267]  = 8'd111;
    TRI_LUT[268]  = 8'd110;
    TRI_LUT[269]  = 8'd109;
    TRI_LUT[270]  = 8'd108;
    TRI_LUT[271]  = 8'd107;
    TRI_LUT[272]  = 8'd106;
    TRI_LUT[273]  = 8'd105;
    TRI_LUT[274]  = 8'd104;
    TRI_LUT[275]  = 8'd103;
    TRI_LUT[276]  = 8'd102;
    TRI_LUT[277]  = 8'd101;
    TRI_LUT[278]  = 8'd100;
    TRI_LUT[279]  = 8'd99;
    TRI_LUT[280]  = 8'd98;
    TRI_LUT[281]  = 8'd97;
    TRI_LUT[282]  = 8'd96;
    TRI_LUT[283]  = 8'd95;
    TRI_LUT[284]  = 8'd94;
    TRI_LUT[285]  = 8'd93;
    TRI_LUT[286]  = 8'd92;
    TRI_LUT[287]  = 8'd91;
    TRI_LUT[288]  = 8'd90;
    TRI_LUT[289]  = 8'd89;
    TRI_LUT[290]  = 8'd88;
    TRI_LUT[291]  = 8'd87;
    TRI_LUT[292]  = 8'd86;
    TRI_LUT[293]  = 8'd85;
    TRI_LUT[294]  = 8'd84;
    TRI_LUT[295]  = 8'd83;
    TRI_LUT[296]  = 8'd82;
    TRI_LUT[297]  = 8'd81;
    TRI_LUT[298]  = 8'd80;
    TRI_LUT[299]  = 8'd79;
    TRI_LUT[300]  = 8'd78;
    TRI_LUT[301]  = 8'd77;
    TRI_LUT[302]  = 8'd76;
    TRI_LUT[303]  = 8'd75;
    TRI_LUT[304]  = 8'd74;
    TRI_LUT[305]  = 8'd73;
    TRI_LUT[306]  = 8'd72;
    TRI_LUT[307]  = 8'd71;
    TRI_LUT[308]  = 8'd70;
    TRI_LUT[309]  = 8'd69;
    TRI_LUT[310]  = 8'd68;
    TRI_LUT[311]  = 8'd67;
    TRI_LUT[312]  = 8'd66;
    TRI_LUT[313]  = 8'd65;
    TRI_LUT[314]  = 8'd64;
    TRI_LUT[315]  = 8'd63;
    TRI_LUT[316]  = 8'd62;
    TRI_LUT[317]  = 8'd61;
    TRI_LUT[318]  = 8'd60;
    TRI_LUT[319]  = 8'd59;
    TRI_LUT[320]  = 8'd58;
    TRI_LUT[321]  = 8'd57;
    TRI_LUT[322]  = 8'd56;
    TRI_LUT[323]  = 8'd54;
    TRI_LUT[324]  = 8'd53;
    TRI_LUT[325]  = 8'd52;
    TRI_LUT[326]  = 8'd51;
    TRI_LUT[327]  = 8'd50;
    TRI_LUT[328]  = 8'd49;
    TRI_LUT[329]  = 8'd48;
    TRI_LUT[330]  = 8'd47;
    TRI_LUT[331]  = 8'd46;
    TRI_LUT[332]  = 8'd45;
    TRI_LUT[333]  = 8'd44;
    TRI_LUT[334]  = 8'd43;
    TRI_LUT[335]  = 8'd42;
    TRI_LUT[336]  = 8'd41;
    TRI_LUT[337]  = 8'd40;
    TRI_LUT[338]  = 8'd39;
    TRI_LUT[339]  = 8'd38;
    TRI_LUT[340]  = 8'd37;
    TRI_LUT[341]  = 8'd36;
    TRI_LUT[342]  = 8'd35;
    TRI_LUT[343]  = 8'd34;
    TRI_LUT[344]  = 8'd33;
    TRI_LUT[345]  = 8'd32;
    TRI_LUT[346]  = 8'd31;
    TRI_LUT[347]  = 8'd30;
    TRI_LUT[348]  = 8'd29;
    TRI_LUT[349]  = 8'd28;
    TRI_LUT[350]  = 8'd27;
    TRI_LUT[351]  = 8'd26;
    TRI_LUT[352]  = 8'd25;
    TRI_LUT[353]  = 8'd24;
    TRI_LUT[354]  = 8'd23;
    TRI_LUT[355]  = 8'd22;
    TRI_LUT[356]  = 8'd21;
    TRI_LUT[357]  = 8'd20;
    TRI_LUT[358]  = 8'd19;
    TRI_LUT[359]  = 8'd18;
    TRI_LUT[360]  = 8'd17;
    TRI_LUT[361]  = 8'd16;
    TRI_LUT[362]  = 8'd15;
    TRI_LUT[363]  = 8'd14;
    TRI_LUT[364]  = 8'd13;
    TRI_LUT[365]  = 8'd12;
    TRI_LUT[366]  = 8'd11;
    TRI_LUT[367]  = 8'd10;
    TRI_LUT[368]  = 8'd9;
    TRI_LUT[369]  = 8'd8;
    TRI_LUT[370]  = 8'd7;
    TRI_LUT[371]  = 8'd6;
    TRI_LUT[372]  = 8'd5;
    TRI_LUT[373]  = 8'd4;
    TRI_LUT[374]  = 8'd3;
    TRI_LUT[375]  = 8'd2;
    TRI_LUT[376]  = 8'd0;
    TRI_LUT[377]  = 8'd1;
    TRI_LUT[378]  = 8'd2;
    TRI_LUT[379]  = 8'd3;
    TRI_LUT[380]  = 8'd4;
    TRI_LUT[381]  = 8'd5;
    TRI_LUT[382]  = 8'd6;
    TRI_LUT[383]  = 8'd7;
    TRI_LUT[384]  = 8'd8;
    TRI_LUT[385]  = 8'd9;
    TRI_LUT[386]  = 8'd10;
    TRI_LUT[387]  = 8'd11;
    TRI_LUT[388]  = 8'd12;
    TRI_LUT[389]  = 8'd13;
    TRI_LUT[390]  = 8'd14;
    TRI_LUT[391]  = 8'd15;
    TRI_LUT[392]  = 8'd16;
    TRI_LUT[393]  = 8'd17;
    TRI_LUT[394]  = 8'd19;
    TRI_LUT[395]  = 8'd20;
    TRI_LUT[396]  = 8'd21;
    TRI_LUT[397]  = 8'd22;
    TRI_LUT[398]  = 8'd23;
    TRI_LUT[399]  = 8'd24;
    TRI_LUT[400]  = 8'd25;
    TRI_LUT[401]  = 8'd26;
    TRI_LUT[402]  = 8'd27;
    TRI_LUT[403]  = 8'd28;
    TRI_LUT[404]  = 8'd29;
    TRI_LUT[405]  = 8'd30;
    TRI_LUT[406]  = 8'd31;
    TRI_LUT[407]  = 8'd32;
    TRI_LUT[408]  = 8'd33;
    TRI_LUT[409]  = 8'd34;
    TRI_LUT[410]  = 8'd35;
    TRI_LUT[411]  = 8'd36;
    TRI_LUT[412]  = 8'd37;
    TRI_LUT[413]  = 8'd38;
    TRI_LUT[414]  = 8'd39;
    TRI_LUT[415]  = 8'd40;
    TRI_LUT[416]  = 8'd41;
    TRI_LUT[417]  = 8'd42;
    TRI_LUT[418]  = 8'd43;
    TRI_LUT[419]  = 8'd44;
    TRI_LUT[420]  = 8'd45;
    TRI_LUT[421]  = 8'd46;
    TRI_LUT[422]  = 8'd47;
    TRI_LUT[423]  = 8'd48;
    TRI_LUT[424]  = 8'd49;
    TRI_LUT[425]  = 8'd50;
    TRI_LUT[426]  = 8'd51;
    TRI_LUT[427]  = 8'd52;
    TRI_LUT[428]  = 8'd53;
    TRI_LUT[429]  = 8'd54;
    TRI_LUT[430]  = 8'd55;
    TRI_LUT[431]  = 8'd56;
    TRI_LUT[432]  = 8'd57;
    TRI_LUT[433]  = 8'd58;
    TRI_LUT[434]  = 8'd59;
    TRI_LUT[435]  = 8'd60;
    TRI_LUT[436]  = 8'd61;
    TRI_LUT[437]  = 8'd62;
    TRI_LUT[438]  = 8'd63;
    TRI_LUT[439]  = 8'd64;
    TRI_LUT[440]  = 8'd65;
    TRI_LUT[441]  = 8'd66;
    TRI_LUT[442]  = 8'd67;
    TRI_LUT[443]  = 8'd68;
    TRI_LUT[444]  = 8'd69;
    TRI_LUT[445]  = 8'd70;
    TRI_LUT[446]  = 8'd71;
    TRI_LUT[447]  = 8'd72;
    TRI_LUT[448]  = 8'd73;
    TRI_LUT[449]  = 8'd74;
    TRI_LUT[450]  = 8'd75;
    TRI_LUT[451]  = 8'd76;
    TRI_LUT[452]  = 8'd77;
    TRI_LUT[453]  = 8'd78;
    TRI_LUT[454]  = 8'd79;
    TRI_LUT[455]  = 8'd80;
    TRI_LUT[456]  = 8'd81;
    TRI_LUT[457]  = 8'd82;
    TRI_LUT[458]  = 8'd83;
    TRI_LUT[459]  = 8'd84;
    TRI_LUT[460]  = 8'd85;
    TRI_LUT[461]  = 8'd86;
    TRI_LUT[462]  = 8'd87;
    TRI_LUT[463]  = 8'd88;
    TRI_LUT[464]  = 8'd89;
    TRI_LUT[465]  = 8'd90;
    TRI_LUT[466]  = 8'd92;
    TRI_LUT[467]  = 8'd93;
    TRI_LUT[468]  = 8'd94;
    TRI_LUT[469]  = 8'd95;
    TRI_LUT[470]  = 8'd96;
    TRI_LUT[471]  = 8'd97;
    TRI_LUT[472]  = 8'd98;
    TRI_LUT[473]  = 8'd99;
    TRI_LUT[474]  = 8'd100;
    TRI_LUT[475]  = 8'd101;
    TRI_LUT[476]  = 8'd102;
    TRI_LUT[477]  = 8'd103;
    TRI_LUT[478]  = 8'd104;
    TRI_LUT[479]  = 8'd105;
    TRI_LUT[480]  = 8'd106;
    TRI_LUT[481]  = 8'd107;
    TRI_LUT[482]  = 8'd108;
    TRI_LUT[483]  = 8'd109;
    TRI_LUT[484]  = 8'd110;
    TRI_LUT[485]  = 8'd111;
    TRI_LUT[486]  = 8'd112;
    TRI_LUT[487]  = 8'd113;
    TRI_LUT[488]  = 8'd114;
    TRI_LUT[489]  = 8'd115;
    TRI_LUT[490]  = 8'd116;
    TRI_LUT[491]  = 8'd117;
    TRI_LUT[492]  = 8'd118;
    TRI_LUT[493]  = 8'd119;
    TRI_LUT[494]  = 8'd120;
    TRI_LUT[495]  = 8'd121;
    TRI_LUT[496]  = 8'd122;
    TRI_LUT[497]  = 8'd123;
    TRI_LUT[498]  = 8'd124;
    TRI_LUT[499]  = 8'd125;
    TRI_LUT[500]  = 8'd126;
end

    
      always_ff @(posedge clk or posedge rst) begin
        if (rst)
          ptr <= 9'd0;
        else if (in_valid) begin
          // compute next pointer, with wrap at MAX_INDEX+1
          nxt = ptr + 9'd1;
          if (nxt > 500)
            ptr <= nxt - 501;
          else
            ptr <= nxt;
        end
      end
   
    // ----------------------------------------------------------------
    // Runtime lookup
    // ----------------------------------------------------------------
    assign out_data = TRI_LUT[ptr];

endmodule
